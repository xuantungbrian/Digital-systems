module DDS();

endmodule