module FFXII_LB_Cursor(RGB,YX);

output reg [11:0]RGB;
input wire [19:0]YX;
parameter Y0X0={10'd0, 10'd0};
parameter Y0X1={10'd0, 10'd1};
parameter Y0X2={10'd0, 10'd2};
parameter Y0X3={10'd0, 10'd3};
parameter Y0X4={10'd0, 10'd4};
parameter Y0X5={10'd0, 10'd5};
parameter Y0X6={10'd0, 10'd6};
parameter Y0X7={10'd0, 10'd7};
parameter Y0X8={10'd0, 10'd8};
parameter Y0X9={10'd0, 10'd9};
parameter Y0X10={10'd0, 10'd10};
parameter Y0X11={10'd0, 10'd11};
parameter Y0X12={10'd0, 10'd12};
parameter Y0X13={10'd0, 10'd13};
parameter Y0X14={10'd0, 10'd14};
parameter Y0X15={10'd0, 10'd15};
parameter Y0X16={10'd0, 10'd16};
parameter Y0X17={10'd0, 10'd17};
parameter Y0X18={10'd0, 10'd18};
parameter Y0X19={10'd0, 10'd19};
parameter Y0X20={10'd0, 10'd20};
parameter Y0X21={10'd0, 10'd21};
parameter Y0X22={10'd0, 10'd22};
parameter Y0X23={10'd0, 10'd23};
parameter Y0X24={10'd0, 10'd24};
parameter Y0X25={10'd0, 10'd25};
parameter Y0X26={10'd0, 10'd26};
parameter Y0X27={10'd0, 10'd27};
parameter Y0X28={10'd0, 10'd28};
parameter Y1X1={10'd1, 10'd1};
parameter Y1X2={10'd1, 10'd2};
parameter Y1X3={10'd1, 10'd3};
parameter Y1X4={10'd1, 10'd4};
parameter Y1X5={10'd1, 10'd5};
parameter Y1X6={10'd1, 10'd6};
parameter Y1X7={10'd1, 10'd7};
parameter Y1X8={10'd1, 10'd8};
parameter Y1X9={10'd1, 10'd9};
parameter Y1X10={10'd1, 10'd10};
parameter Y1X11={10'd1, 10'd11};
parameter Y1X12={10'd1, 10'd12};
parameter Y1X13={10'd1, 10'd13};
parameter Y1X14={10'd1, 10'd14};
parameter Y1X15={10'd1, 10'd15};
parameter Y1X16={10'd1, 10'd16};
parameter Y1X17={10'd1, 10'd17};
parameter Y1X18={10'd1, 10'd18};
parameter Y1X19={10'd1, 10'd19};
parameter Y1X20={10'd1, 10'd20};
parameter Y1X21={10'd1, 10'd21};
parameter Y1X22={10'd1, 10'd22};
parameter Y1X23={10'd1, 10'd23};
parameter Y1X24={10'd1, 10'd24};
parameter Y1X25={10'd1, 10'd25};
parameter Y1X26={10'd1, 10'd26};
parameter Y1X27={10'd1, 10'd27};
parameter Y1X28={10'd1, 10'd28};
parameter Y2X1={10'd2, 10'd1};
parameter Y2X2={10'd2, 10'd2};
parameter Y2X3={10'd2, 10'd3};
parameter Y2X4={10'd2, 10'd4};
parameter Y2X5={10'd2, 10'd5};
parameter Y2X6={10'd2, 10'd6};
parameter Y2X7={10'd2, 10'd7};
parameter Y2X8={10'd2, 10'd8};
parameter Y2X9={10'd2, 10'd9};
parameter Y2X10={10'd2, 10'd10};
parameter Y2X11={10'd2, 10'd11};
parameter Y2X12={10'd2, 10'd12};
parameter Y2X13={10'd2, 10'd13};
parameter Y2X14={10'd2, 10'd14};
parameter Y2X15={10'd2, 10'd15};
parameter Y2X16={10'd2, 10'd16};
parameter Y2X17={10'd2, 10'd17};
parameter Y2X18={10'd2, 10'd18};
parameter Y2X19={10'd2, 10'd19};
parameter Y2X20={10'd2, 10'd20};
parameter Y2X21={10'd2, 10'd21};
parameter Y2X22={10'd2, 10'd22};
parameter Y2X23={10'd2, 10'd23};
parameter Y2X24={10'd2, 10'd24};
parameter Y2X25={10'd2, 10'd25};
parameter Y2X26={10'd2, 10'd26};
parameter Y2X27={10'd2, 10'd27};
parameter Y2X28={10'd2, 10'd28};
parameter Y3X1={10'd3, 10'd1};
parameter Y3X2={10'd3, 10'd2};
parameter Y3X3={10'd3, 10'd3};
parameter Y3X4={10'd3, 10'd4};
parameter Y3X5={10'd3, 10'd5};
parameter Y3X6={10'd3, 10'd6};
parameter Y3X7={10'd3, 10'd7};
parameter Y3X8={10'd3, 10'd8};
parameter Y3X9={10'd3, 10'd9};
parameter Y3X10={10'd3, 10'd10};
parameter Y3X11={10'd3, 10'd11};
parameter Y3X12={10'd3, 10'd12};
parameter Y3X13={10'd3, 10'd13};
parameter Y3X14={10'd3, 10'd14};
parameter Y3X15={10'd3, 10'd15};
parameter Y3X16={10'd3, 10'd16};
parameter Y3X17={10'd3, 10'd17};
parameter Y3X18={10'd3, 10'd18};
parameter Y3X19={10'd3, 10'd19};
parameter Y3X20={10'd3, 10'd20};
parameter Y3X21={10'd3, 10'd21};
parameter Y3X22={10'd3, 10'd22};
parameter Y3X23={10'd3, 10'd23};
parameter Y3X24={10'd3, 10'd24};
parameter Y3X25={10'd3, 10'd25};
parameter Y3X26={10'd3, 10'd26};
parameter Y3X27={10'd3, 10'd27};
parameter Y3X28={10'd3, 10'd28};
parameter Y4X1={10'd4, 10'd1};
parameter Y4X2={10'd4, 10'd2};
parameter Y4X3={10'd4, 10'd3};
parameter Y4X4={10'd4, 10'd4};
parameter Y4X5={10'd4, 10'd5};
parameter Y4X6={10'd4, 10'd6};
parameter Y4X7={10'd4, 10'd7};
parameter Y4X8={10'd4, 10'd8};
parameter Y4X9={10'd4, 10'd9};
parameter Y4X10={10'd4, 10'd10};
parameter Y4X11={10'd4, 10'd11};
parameter Y4X12={10'd4, 10'd12};
parameter Y4X13={10'd4, 10'd13};
parameter Y4X14={10'd4, 10'd14};
parameter Y4X15={10'd4, 10'd15};
parameter Y4X16={10'd4, 10'd16};
parameter Y4X17={10'd4, 10'd17};
parameter Y4X18={10'd4, 10'd18};
parameter Y4X19={10'd4, 10'd19};
parameter Y4X20={10'd4, 10'd20};
parameter Y4X21={10'd4, 10'd21};
parameter Y4X22={10'd4, 10'd22};
parameter Y4X23={10'd4, 10'd23};
parameter Y4X24={10'd4, 10'd24};
parameter Y4X25={10'd4, 10'd25};
parameter Y4X26={10'd4, 10'd26};
parameter Y4X27={10'd4, 10'd27};
parameter Y4X28={10'd4, 10'd28};
parameter Y5X1={10'd5, 10'd1};
parameter Y5X2={10'd5, 10'd2};
parameter Y5X3={10'd5, 10'd3};
parameter Y5X4={10'd5, 10'd4};
parameter Y5X5={10'd5, 10'd5};
parameter Y5X6={10'd5, 10'd6};
parameter Y5X7={10'd5, 10'd7};
parameter Y5X8={10'd5, 10'd8};
parameter Y5X9={10'd5, 10'd9};
parameter Y5X10={10'd5, 10'd10};
parameter Y5X11={10'd5, 10'd11};
parameter Y5X12={10'd5, 10'd12};
parameter Y5X13={10'd5, 10'd13};
parameter Y5X14={10'd5, 10'd14};
parameter Y5X15={10'd5, 10'd15};
parameter Y5X16={10'd5, 10'd16};
parameter Y5X17={10'd5, 10'd17};
parameter Y5X18={10'd5, 10'd18};
parameter Y5X19={10'd5, 10'd19};
parameter Y5X20={10'd5, 10'd20};
parameter Y5X21={10'd5, 10'd21};
parameter Y5X22={10'd5, 10'd22};
parameter Y5X23={10'd5, 10'd23};
parameter Y5X24={10'd5, 10'd24};
parameter Y5X25={10'd5, 10'd25};
parameter Y5X26={10'd5, 10'd26};
parameter Y5X27={10'd5, 10'd27};
parameter Y5X28={10'd5, 10'd28};
parameter Y6X1={10'd6, 10'd1};
parameter Y6X2={10'd6, 10'd2};
parameter Y6X3={10'd6, 10'd3};
parameter Y6X4={10'd6, 10'd4};
parameter Y6X5={10'd6, 10'd5};
parameter Y6X6={10'd6, 10'd6};
parameter Y6X7={10'd6, 10'd7};
parameter Y6X8={10'd6, 10'd8};
parameter Y6X9={10'd6, 10'd9};
parameter Y6X10={10'd6, 10'd10};
parameter Y6X11={10'd6, 10'd11};
parameter Y6X12={10'd6, 10'd12};
parameter Y6X13={10'd6, 10'd13};
parameter Y6X14={10'd6, 10'd14};
parameter Y6X15={10'd6, 10'd15};
parameter Y6X16={10'd6, 10'd16};
parameter Y6X17={10'd6, 10'd17};
parameter Y6X18={10'd6, 10'd18};
parameter Y6X19={10'd6, 10'd19};
parameter Y6X20={10'd6, 10'd20};
parameter Y6X21={10'd6, 10'd21};
parameter Y6X22={10'd6, 10'd22};
parameter Y6X23={10'd6, 10'd23};
parameter Y6X24={10'd6, 10'd24};
parameter Y6X25={10'd6, 10'd25};
parameter Y6X26={10'd6, 10'd26};
parameter Y6X27={10'd6, 10'd27};
parameter Y6X28={10'd6, 10'd28};
parameter Y7X1={10'd7, 10'd1};
parameter Y7X2={10'd7, 10'd2};
parameter Y7X3={10'd7, 10'd3};
parameter Y7X4={10'd7, 10'd4};
parameter Y7X5={10'd7, 10'd5};
parameter Y7X6={10'd7, 10'd6};
parameter Y7X7={10'd7, 10'd7};
parameter Y7X8={10'd7, 10'd8};
parameter Y7X9={10'd7, 10'd9};
parameter Y7X10={10'd7, 10'd10};
parameter Y7X11={10'd7, 10'd11};
parameter Y7X12={10'd7, 10'd12};
parameter Y7X13={10'd7, 10'd13};
parameter Y7X14={10'd7, 10'd14};
parameter Y7X15={10'd7, 10'd15};
parameter Y7X16={10'd7, 10'd16};
parameter Y7X17={10'd7, 10'd17};
parameter Y7X18={10'd7, 10'd18};
parameter Y7X19={10'd7, 10'd19};
parameter Y7X20={10'd7, 10'd20};
parameter Y7X21={10'd7, 10'd21};
parameter Y7X22={10'd7, 10'd22};
parameter Y7X23={10'd7, 10'd23};
parameter Y7X24={10'd7, 10'd24};
parameter Y7X25={10'd7, 10'd25};
parameter Y7X26={10'd7, 10'd26};
parameter Y7X27={10'd7, 10'd27};
parameter Y7X28={10'd7, 10'd28};
parameter Y8X1={10'd8, 10'd1};
parameter Y8X2={10'd8, 10'd2};
parameter Y8X3={10'd8, 10'd3};
parameter Y8X4={10'd8, 10'd4};
parameter Y8X5={10'd8, 10'd5};
parameter Y8X6={10'd8, 10'd6};
parameter Y8X7={10'd8, 10'd7};
parameter Y8X8={10'd8, 10'd8};
parameter Y8X9={10'd8, 10'd9};
parameter Y8X10={10'd8, 10'd10};
parameter Y8X11={10'd8, 10'd11};
parameter Y8X12={10'd8, 10'd12};
parameter Y8X13={10'd8, 10'd13};
parameter Y8X14={10'd8, 10'd14};
parameter Y8X15={10'd8, 10'd15};
parameter Y8X16={10'd8, 10'd16};
parameter Y8X17={10'd8, 10'd17};
parameter Y8X18={10'd8, 10'd18};
parameter Y8X19={10'd8, 10'd19};
parameter Y8X20={10'd8, 10'd20};
parameter Y8X21={10'd8, 10'd21};
parameter Y8X22={10'd8, 10'd22};
parameter Y8X23={10'd8, 10'd23};
parameter Y8X24={10'd8, 10'd24};
parameter Y8X25={10'd8, 10'd25};
parameter Y8X26={10'd8, 10'd26};
parameter Y8X27={10'd8, 10'd27};
parameter Y8X28={10'd8, 10'd28};
parameter Y9X1={10'd9, 10'd1};
parameter Y9X2={10'd9, 10'd2};
parameter Y9X3={10'd9, 10'd3};
parameter Y9X4={10'd9, 10'd4};
parameter Y9X5={10'd9, 10'd5};
parameter Y9X6={10'd9, 10'd6};
parameter Y9X7={10'd9, 10'd7};
parameter Y9X8={10'd9, 10'd8};
parameter Y9X9={10'd9, 10'd9};
parameter Y9X10={10'd9, 10'd10};
parameter Y9X11={10'd9, 10'd11};
parameter Y9X12={10'd9, 10'd12};
parameter Y9X13={10'd9, 10'd13};
parameter Y9X14={10'd9, 10'd14};
parameter Y9X15={10'd9, 10'd15};
parameter Y9X16={10'd9, 10'd16};
parameter Y9X17={10'd9, 10'd17};
parameter Y9X18={10'd9, 10'd18};
parameter Y9X19={10'd9, 10'd19};
parameter Y9X20={10'd9, 10'd20};
parameter Y9X21={10'd9, 10'd21};
parameter Y9X22={10'd9, 10'd22};
parameter Y9X23={10'd9, 10'd23};
parameter Y9X24={10'd9, 10'd24};
parameter Y9X25={10'd9, 10'd25};
parameter Y9X26={10'd9, 10'd26};
parameter Y9X27={10'd9, 10'd27};
parameter Y9X28={10'd9, 10'd28};
parameter Y10X1={10'd10, 10'd1};
parameter Y10X2={10'd10, 10'd2};
parameter Y10X3={10'd10, 10'd3};
parameter Y10X4={10'd10, 10'd4};
parameter Y10X5={10'd10, 10'd5};
parameter Y10X6={10'd10, 10'd6};
parameter Y10X7={10'd10, 10'd7};
parameter Y10X8={10'd10, 10'd8};
parameter Y10X9={10'd10, 10'd9};
parameter Y10X10={10'd10, 10'd10};
parameter Y10X11={10'd10, 10'd11};
parameter Y10X12={10'd10, 10'd12};
parameter Y10X13={10'd10, 10'd13};
parameter Y10X14={10'd10, 10'd14};
parameter Y10X15={10'd10, 10'd15};
parameter Y10X16={10'd10, 10'd16};
parameter Y10X17={10'd10, 10'd17};
parameter Y10X18={10'd10, 10'd18};
parameter Y10X19={10'd10, 10'd19};
parameter Y10X20={10'd10, 10'd20};
parameter Y10X21={10'd10, 10'd21};
parameter Y10X22={10'd10, 10'd22};
parameter Y10X23={10'd10, 10'd23};
parameter Y10X24={10'd10, 10'd24};
parameter Y10X25={10'd10, 10'd25};
parameter Y10X26={10'd10, 10'd26};
parameter Y10X27={10'd10, 10'd27};
parameter Y10X28={10'd10, 10'd28};
parameter Y11X1={10'd11, 10'd1};
parameter Y11X2={10'd11, 10'd2};
parameter Y11X3={10'd11, 10'd3};
parameter Y11X4={10'd11, 10'd4};
parameter Y11X5={10'd11, 10'd5};
parameter Y11X6={10'd11, 10'd6};
parameter Y11X7={10'd11, 10'd7};
parameter Y11X8={10'd11, 10'd8};
parameter Y11X9={10'd11, 10'd9};
parameter Y11X10={10'd11, 10'd10};
parameter Y11X11={10'd11, 10'd11};
parameter Y11X12={10'd11, 10'd12};
parameter Y11X13={10'd11, 10'd13};
parameter Y11X14={10'd11, 10'd14};
parameter Y11X15={10'd11, 10'd15};
parameter Y11X16={10'd11, 10'd16};
parameter Y11X17={10'd11, 10'd17};
parameter Y11X18={10'd11, 10'd18};
parameter Y11X19={10'd11, 10'd19};
parameter Y11X20={10'd11, 10'd20};
parameter Y11X21={10'd11, 10'd21};
parameter Y11X22={10'd11, 10'd22};
parameter Y11X23={10'd11, 10'd23};
parameter Y11X24={10'd11, 10'd24};
parameter Y11X25={10'd11, 10'd25};
parameter Y11X26={10'd11, 10'd26};
parameter Y11X27={10'd11, 10'd27};
parameter Y11X28={10'd11, 10'd28};
parameter Y12X1={10'd12, 10'd1};
parameter Y12X2={10'd12, 10'd2};
parameter Y12X3={10'd12, 10'd3};
parameter Y12X4={10'd12, 10'd4};
parameter Y12X5={10'd12, 10'd5};
parameter Y12X6={10'd12, 10'd6};
parameter Y12X7={10'd12, 10'd7};
parameter Y12X8={10'd12, 10'd8};
parameter Y12X9={10'd12, 10'd9};
parameter Y12X10={10'd12, 10'd10};
parameter Y12X11={10'd12, 10'd11};
parameter Y12X12={10'd12, 10'd12};
parameter Y12X13={10'd12, 10'd13};
parameter Y12X14={10'd12, 10'd14};
parameter Y12X15={10'd12, 10'd15};
parameter Y12X16={10'd12, 10'd16};
parameter Y12X17={10'd12, 10'd17};
parameter Y12X18={10'd12, 10'd18};
parameter Y12X19={10'd12, 10'd19};
parameter Y12X20={10'd12, 10'd20};
parameter Y12X21={10'd12, 10'd21};
parameter Y12X22={10'd12, 10'd22};
parameter Y12X23={10'd12, 10'd23};
parameter Y12X24={10'd12, 10'd24};
parameter Y12X25={10'd12, 10'd25};
parameter Y12X26={10'd12, 10'd26};
parameter Y12X27={10'd12, 10'd27};
parameter Y12X28={10'd12, 10'd28};
parameter Y13X1={10'd13, 10'd1};
parameter Y13X2={10'd13, 10'd2};
parameter Y13X3={10'd13, 10'd3};
parameter Y13X4={10'd13, 10'd4};
parameter Y13X5={10'd13, 10'd5};
parameter Y13X6={10'd13, 10'd6};
parameter Y13X7={10'd13, 10'd7};
parameter Y13X8={10'd13, 10'd8};
parameter Y13X9={10'd13, 10'd9};
parameter Y13X10={10'd13, 10'd10};
parameter Y13X11={10'd13, 10'd11};
parameter Y13X12={10'd13, 10'd12};
parameter Y13X13={10'd13, 10'd13};
parameter Y13X14={10'd13, 10'd14};
parameter Y13X15={10'd13, 10'd15};
parameter Y13X16={10'd13, 10'd16};
parameter Y13X17={10'd13, 10'd17};
parameter Y13X18={10'd13, 10'd18};
parameter Y13X19={10'd13, 10'd19};
parameter Y13X20={10'd13, 10'd20};
parameter Y13X21={10'd13, 10'd21};
parameter Y13X22={10'd13, 10'd22};
parameter Y13X23={10'd13, 10'd23};
parameter Y13X24={10'd13, 10'd24};
parameter Y13X25={10'd13, 10'd25};
parameter Y13X26={10'd13, 10'd26};
parameter Y13X27={10'd13, 10'd27};
parameter Y13X28={10'd13, 10'd28};
parameter Y14X1={10'd14, 10'd1};
parameter Y14X2={10'd14, 10'd2};
parameter Y14X3={10'd14, 10'd3};
parameter Y14X4={10'd14, 10'd4};
parameter Y14X5={10'd14, 10'd5};
parameter Y14X6={10'd14, 10'd6};
parameter Y14X7={10'd14, 10'd7};
parameter Y14X8={10'd14, 10'd8};
parameter Y14X9={10'd14, 10'd9};
parameter Y14X10={10'd14, 10'd10};
parameter Y14X11={10'd14, 10'd11};
parameter Y14X12={10'd14, 10'd12};
parameter Y14X13={10'd14, 10'd13};
parameter Y14X14={10'd14, 10'd14};
parameter Y14X15={10'd14, 10'd15};
parameter Y14X16={10'd14, 10'd16};
parameter Y14X17={10'd14, 10'd17};
parameter Y14X18={10'd14, 10'd18};
parameter Y14X19={10'd14, 10'd19};
parameter Y14X20={10'd14, 10'd20};
parameter Y14X21={10'd14, 10'd21};
parameter Y14X22={10'd14, 10'd22};
parameter Y14X23={10'd14, 10'd23};
parameter Y14X24={10'd14, 10'd24};
parameter Y14X25={10'd14, 10'd25};
parameter Y14X26={10'd14, 10'd26};
parameter Y14X27={10'd14, 10'd27};
parameter Y14X28={10'd14, 10'd28};
parameter Y15X1={10'd15, 10'd1};
parameter Y15X2={10'd15, 10'd2};
parameter Y15X3={10'd15, 10'd3};
parameter Y15X4={10'd15, 10'd4};
parameter Y15X5={10'd15, 10'd5};
parameter Y15X6={10'd15, 10'd6};
parameter Y15X7={10'd15, 10'd7};
parameter Y15X8={10'd15, 10'd8};
parameter Y15X9={10'd15, 10'd9};
parameter Y15X10={10'd15, 10'd10};
parameter Y15X11={10'd15, 10'd11};
parameter Y15X12={10'd15, 10'd12};
parameter Y15X13={10'd15, 10'd13};
parameter Y15X14={10'd15, 10'd14};
parameter Y15X15={10'd15, 10'd15};
parameter Y15X16={10'd15, 10'd16};
parameter Y15X17={10'd15, 10'd17};
parameter Y15X18={10'd15, 10'd18};
parameter Y15X19={10'd15, 10'd19};
parameter Y15X20={10'd15, 10'd20};
parameter Y15X21={10'd15, 10'd21};
parameter Y15X22={10'd15, 10'd22};
parameter Y15X23={10'd15, 10'd23};
parameter Y15X24={10'd15, 10'd24};
parameter Y15X25={10'd15, 10'd25};
parameter Y15X26={10'd15, 10'd26};
parameter Y15X27={10'd15, 10'd27};
parameter Y15X28={10'd15, 10'd28};
parameter Y16X1={10'd16, 10'd1};
parameter Y16X2={10'd16, 10'd2};
parameter Y16X3={10'd16, 10'd3};
parameter Y16X4={10'd16, 10'd4};
parameter Y16X5={10'd16, 10'd5};
parameter Y16X6={10'd16, 10'd6};
parameter Y16X7={10'd16, 10'd7};
parameter Y16X8={10'd16, 10'd8};
parameter Y16X9={10'd16, 10'd9};
parameter Y16X10={10'd16, 10'd10};
parameter Y16X11={10'd16, 10'd11};
parameter Y16X12={10'd16, 10'd12};
parameter Y16X13={10'd16, 10'd13};
parameter Y16X14={10'd16, 10'd14};
parameter Y16X15={10'd16, 10'd15};
parameter Y16X16={10'd16, 10'd16};
parameter Y16X17={10'd16, 10'd17};
parameter Y16X18={10'd16, 10'd18};
parameter Y16X19={10'd16, 10'd19};
parameter Y16X20={10'd16, 10'd20};
parameter Y16X21={10'd16, 10'd21};
parameter Y16X22={10'd16, 10'd22};
parameter Y16X23={10'd16, 10'd23};
parameter Y16X24={10'd16, 10'd24};
parameter Y16X25={10'd16, 10'd25};
parameter Y16X26={10'd16, 10'd26};
parameter Y16X27={10'd16, 10'd27};
parameter Y16X28={10'd16, 10'd28};
parameter Y17X1={10'd17, 10'd1};
parameter Y17X2={10'd17, 10'd2};
parameter Y17X3={10'd17, 10'd3};
parameter Y17X4={10'd17, 10'd4};
parameter Y17X5={10'd17, 10'd5};
parameter Y17X6={10'd17, 10'd6};
parameter Y17X7={10'd17, 10'd7};
parameter Y17X8={10'd17, 10'd8};
parameter Y17X9={10'd17, 10'd9};
parameter Y17X10={10'd17, 10'd10};
parameter Y17X11={10'd17, 10'd11};
parameter Y17X12={10'd17, 10'd12};
parameter Y17X13={10'd17, 10'd13};
parameter Y17X14={10'd17, 10'd14};
parameter Y17X15={10'd17, 10'd15};
parameter Y17X16={10'd17, 10'd16};
parameter Y17X17={10'd17, 10'd17};
parameter Y17X18={10'd17, 10'd18};
parameter Y17X19={10'd17, 10'd19};
parameter Y17X20={10'd17, 10'd20};
parameter Y17X21={10'd17, 10'd21};
parameter Y17X22={10'd17, 10'd22};
parameter Y17X23={10'd17, 10'd23};
parameter Y17X24={10'd17, 10'd24};
parameter Y17X25={10'd17, 10'd25};
parameter Y17X26={10'd17, 10'd26};
parameter Y17X27={10'd17, 10'd27};
parameter Y17X28={10'd17, 10'd28};
parameter Y18X1={10'd18, 10'd1};
parameter Y18X2={10'd18, 10'd2};
parameter Y18X3={10'd18, 10'd3};
parameter Y18X4={10'd18, 10'd4};
parameter Y18X5={10'd18, 10'd5};
parameter Y18X6={10'd18, 10'd6};
parameter Y18X7={10'd18, 10'd7};
parameter Y18X8={10'd18, 10'd8};
parameter Y18X9={10'd18, 10'd9};
parameter Y18X10={10'd18, 10'd10};
parameter Y18X11={10'd18, 10'd11};
parameter Y18X12={10'd18, 10'd12};
parameter Y18X13={10'd18, 10'd13};
parameter Y18X14={10'd18, 10'd14};
parameter Y18X15={10'd18, 10'd15};
parameter Y18X16={10'd18, 10'd16};
parameter Y18X17={10'd18, 10'd17};
parameter Y18X18={10'd18, 10'd18};
parameter Y18X19={10'd18, 10'd19};
parameter Y18X20={10'd18, 10'd20};
parameter Y18X21={10'd18, 10'd21};
parameter Y18X22={10'd18, 10'd22};
parameter Y18X23={10'd18, 10'd23};
parameter Y18X24={10'd18, 10'd24};
parameter Y18X25={10'd18, 10'd25};
parameter Y18X26={10'd18, 10'd26};
parameter Y18X27={10'd18, 10'd27};
parameter Y18X28={10'd18, 10'd28};
parameter Y19X1={10'd19, 10'd1};
parameter Y19X2={10'd19, 10'd2};
parameter Y19X3={10'd19, 10'd3};
parameter Y19X4={10'd19, 10'd4};
parameter Y19X5={10'd19, 10'd5};
parameter Y19X6={10'd19, 10'd6};
parameter Y19X7={10'd19, 10'd7};
parameter Y19X8={10'd19, 10'd8};
parameter Y19X9={10'd19, 10'd9};
parameter Y19X10={10'd19, 10'd10};
parameter Y19X11={10'd19, 10'd11};
parameter Y19X12={10'd19, 10'd12};
parameter Y19X13={10'd19, 10'd13};
parameter Y19X14={10'd19, 10'd14};
parameter Y19X15={10'd19, 10'd15};
parameter Y19X16={10'd19, 10'd16};
parameter Y19X17={10'd19, 10'd17};
parameter Y19X18={10'd19, 10'd18};
parameter Y19X19={10'd19, 10'd19};
parameter Y19X20={10'd19, 10'd20};
parameter Y19X21={10'd19, 10'd21};
parameter Y19X22={10'd19, 10'd22};
parameter Y19X23={10'd19, 10'd23};
parameter Y19X24={10'd19, 10'd24};
parameter Y19X25={10'd19, 10'd25};
parameter Y19X26={10'd19, 10'd26};
parameter Y19X27={10'd19, 10'd27};
parameter Y19X28={10'd19, 10'd28};
parameter Y20X1={10'd20, 10'd1};
parameter Y20X2={10'd20, 10'd2};
parameter Y20X3={10'd20, 10'd3};
parameter Y20X4={10'd20, 10'd4};
parameter Y20X5={10'd20, 10'd5};
parameter Y20X6={10'd20, 10'd6};
parameter Y20X7={10'd20, 10'd7};
parameter Y20X8={10'd20, 10'd8};
parameter Y20X9={10'd20, 10'd9};
parameter Y20X10={10'd20, 10'd10};
parameter Y20X11={10'd20, 10'd11};
parameter Y20X12={10'd20, 10'd12};
parameter Y20X13={10'd20, 10'd13};
parameter Y20X14={10'd20, 10'd14};
parameter Y20X15={10'd20, 10'd15};
parameter Y20X16={10'd20, 10'd16};
parameter Y20X17={10'd20, 10'd17};
parameter Y20X18={10'd20, 10'd18};
parameter Y20X19={10'd20, 10'd19};
parameter Y20X20={10'd20, 10'd20};
parameter Y20X21={10'd20, 10'd21};
parameter Y20X22={10'd20, 10'd22};
parameter Y20X23={10'd20, 10'd23};
parameter Y20X24={10'd20, 10'd24};
parameter Y20X25={10'd20, 10'd25};
parameter Y20X26={10'd20, 10'd26};
parameter Y20X27={10'd20, 10'd27};
parameter Y20X28={10'd20, 10'd28};
parameter Y21X1={10'd21, 10'd1};
parameter Y21X2={10'd21, 10'd2};
parameter Y21X3={10'd21, 10'd3};
parameter Y21X4={10'd21, 10'd4};
parameter Y21X5={10'd21, 10'd5};
parameter Y21X6={10'd21, 10'd6};
parameter Y21X7={10'd21, 10'd7};
parameter Y21X8={10'd21, 10'd8};
parameter Y21X9={10'd21, 10'd9};
parameter Y21X10={10'd21, 10'd10};
parameter Y21X11={10'd21, 10'd11};
parameter Y21X12={10'd21, 10'd12};
parameter Y21X13={10'd21, 10'd13};
parameter Y21X14={10'd21, 10'd14};
parameter Y21X15={10'd21, 10'd15};
parameter Y21X16={10'd21, 10'd16};
parameter Y21X17={10'd21, 10'd17};
parameter Y21X18={10'd21, 10'd18};
parameter Y21X19={10'd21, 10'd19};
parameter Y21X20={10'd21, 10'd20};
parameter Y21X21={10'd21, 10'd21};
parameter Y21X22={10'd21, 10'd22};
parameter Y21X23={10'd21, 10'd23};
parameter Y21X24={10'd21, 10'd24};
parameter Y21X25={10'd21, 10'd25};
parameter Y21X26={10'd21, 10'd26};
parameter Y21X27={10'd21, 10'd27};
parameter Y21X28={10'd21, 10'd28};
parameter Y22X1={10'd22, 10'd1};
parameter Y22X2={10'd22, 10'd2};
parameter Y22X3={10'd22, 10'd3};
parameter Y22X4={10'd22, 10'd4};
parameter Y22X5={10'd22, 10'd5};
parameter Y22X6={10'd22, 10'd6};
parameter Y22X7={10'd22, 10'd7};
parameter Y22X8={10'd22, 10'd8};
parameter Y22X9={10'd22, 10'd9};
parameter Y22X10={10'd22, 10'd10};
parameter Y22X11={10'd22, 10'd11};
parameter Y22X12={10'd22, 10'd12};
parameter Y22X13={10'd22, 10'd13};
parameter Y22X14={10'd22, 10'd14};
parameter Y22X15={10'd22, 10'd15};
parameter Y22X16={10'd22, 10'd16};
parameter Y22X17={10'd22, 10'd17};
parameter Y22X18={10'd22, 10'd18};
parameter Y22X19={10'd22, 10'd19};
parameter Y22X20={10'd22, 10'd20};
parameter Y22X21={10'd22, 10'd21};
parameter Y22X22={10'd22, 10'd22};
parameter Y22X23={10'd22, 10'd23};
parameter Y22X24={10'd22, 10'd24};
parameter Y22X25={10'd22, 10'd25};
parameter Y22X26={10'd22, 10'd26};
parameter Y22X27={10'd22, 10'd27};
parameter Y22X28={10'd22, 10'd28};
parameter Y23X1={10'd23, 10'd1};
parameter Y23X2={10'd23, 10'd2};
parameter Y23X3={10'd23, 10'd3};
parameter Y23X4={10'd23, 10'd4};
parameter Y23X5={10'd23, 10'd5};
parameter Y23X6={10'd23, 10'd6};
parameter Y23X7={10'd23, 10'd7};
parameter Y23X8={10'd23, 10'd8};
parameter Y23X9={10'd23, 10'd9};
parameter Y23X10={10'd23, 10'd10};
parameter Y23X11={10'd23, 10'd11};
parameter Y23X12={10'd23, 10'd12};
parameter Y23X13={10'd23, 10'd13};
parameter Y23X14={10'd23, 10'd14};
parameter Y23X15={10'd23, 10'd15};
parameter Y23X16={10'd23, 10'd16};
parameter Y23X17={10'd23, 10'd17};
parameter Y23X18={10'd23, 10'd18};
parameter Y23X19={10'd23, 10'd19};
parameter Y23X20={10'd23, 10'd20};
parameter Y23X21={10'd23, 10'd21};
parameter Y23X22={10'd23, 10'd22};
parameter Y23X23={10'd23, 10'd23};
parameter Y23X24={10'd23, 10'd24};
parameter Y23X25={10'd23, 10'd25};
parameter Y23X26={10'd23, 10'd26};
parameter Y23X27={10'd23, 10'd27};
parameter Y23X28={10'd23, 10'd28};
parameter Y24X1={10'd24, 10'd1};
parameter Y24X2={10'd24, 10'd2};
parameter Y24X3={10'd24, 10'd3};
parameter Y24X4={10'd24, 10'd4};
parameter Y24X5={10'd24, 10'd5};
parameter Y24X6={10'd24, 10'd6};
parameter Y24X7={10'd24, 10'd7};
parameter Y24X8={10'd24, 10'd8};
parameter Y24X9={10'd24, 10'd9};
parameter Y24X10={10'd24, 10'd10};
parameter Y24X11={10'd24, 10'd11};
parameter Y24X12={10'd24, 10'd12};
parameter Y24X13={10'd24, 10'd13};
parameter Y24X14={10'd24, 10'd14};
parameter Y24X15={10'd24, 10'd15};
parameter Y24X16={10'd24, 10'd16};
parameter Y24X17={10'd24, 10'd17};
parameter Y24X18={10'd24, 10'd18};
parameter Y24X19={10'd24, 10'd19};
parameter Y24X20={10'd24, 10'd20};
parameter Y24X21={10'd24, 10'd21};
parameter Y24X22={10'd24, 10'd22};
parameter Y24X23={10'd24, 10'd23};
parameter Y24X24={10'd24, 10'd24};
parameter Y24X25={10'd24, 10'd25};
parameter Y24X26={10'd24, 10'd26};
parameter Y24X27={10'd24, 10'd27};
parameter Y24X28={10'd24, 10'd28};
parameter Y25X1={10'd25, 10'd1};
parameter Y25X2={10'd25, 10'd2};
parameter Y25X3={10'd25, 10'd3};
parameter Y25X4={10'd25, 10'd4};
parameter Y25X5={10'd25, 10'd5};
parameter Y25X6={10'd25, 10'd6};
parameter Y25X7={10'd25, 10'd7};
parameter Y25X8={10'd25, 10'd8};
parameter Y25X9={10'd25, 10'd9};
parameter Y25X10={10'd25, 10'd10};
parameter Y25X11={10'd25, 10'd11};
parameter Y25X12={10'd25, 10'd12};
parameter Y25X13={10'd25, 10'd13};
parameter Y25X14={10'd25, 10'd14};
parameter Y25X15={10'd25, 10'd15};
parameter Y25X16={10'd25, 10'd16};
parameter Y25X17={10'd25, 10'd17};
parameter Y25X18={10'd25, 10'd18};
parameter Y25X19={10'd25, 10'd19};
parameter Y25X20={10'd25, 10'd20};
parameter Y25X21={10'd25, 10'd21};
parameter Y25X22={10'd25, 10'd22};
parameter Y25X23={10'd25, 10'd23};
parameter Y25X24={10'd25, 10'd24};
parameter Y25X25={10'd25, 10'd25};
parameter Y25X26={10'd25, 10'd26};
parameter Y25X27={10'd25, 10'd27};
parameter Y25X28={10'd25, 10'd28};
parameter Y26X1={10'd26, 10'd1};
parameter Y26X2={10'd26, 10'd2};
parameter Y26X3={10'd26, 10'd3};
parameter Y26X4={10'd26, 10'd4};
parameter Y26X5={10'd26, 10'd5};
parameter Y26X6={10'd26, 10'd6};
parameter Y26X7={10'd26, 10'd7};
parameter Y26X8={10'd26, 10'd8};
parameter Y26X9={10'd26, 10'd9};
parameter Y26X10={10'd26, 10'd10};
parameter Y26X11={10'd26, 10'd11};
parameter Y26X12={10'd26, 10'd12};
parameter Y26X13={10'd26, 10'd13};
parameter Y26X14={10'd26, 10'd14};
parameter Y26X15={10'd26, 10'd15};
parameter Y26X16={10'd26, 10'd16};
parameter Y26X17={10'd26, 10'd17};
parameter Y26X18={10'd26, 10'd18};
parameter Y26X19={10'd26, 10'd19};
parameter Y26X20={10'd26, 10'd20};
parameter Y26X21={10'd26, 10'd21};
parameter Y26X22={10'd26, 10'd22};
parameter Y26X23={10'd26, 10'd23};
parameter Y26X24={10'd26, 10'd24};
parameter Y26X25={10'd26, 10'd25};
parameter Y26X26={10'd26, 10'd26};
parameter Y26X27={10'd26, 10'd27};
parameter Y26X28={10'd26, 10'd28};
parameter Y27X1={10'd27, 10'd1};
parameter Y27X2={10'd27, 10'd2};
parameter Y27X3={10'd27, 10'd3};
parameter Y27X4={10'd27, 10'd4};
parameter Y27X5={10'd27, 10'd5};
parameter Y27X6={10'd27, 10'd6};
parameter Y27X7={10'd27, 10'd7};
parameter Y27X8={10'd27, 10'd8};
parameter Y27X9={10'd27, 10'd9};
parameter Y27X10={10'd27, 10'd10};
parameter Y27X11={10'd27, 10'd11};
parameter Y27X12={10'd27, 10'd12};
parameter Y27X13={10'd27, 10'd13};
parameter Y27X14={10'd27, 10'd14};
parameter Y27X15={10'd27, 10'd15};
parameter Y27X16={10'd27, 10'd16};
parameter Y27X17={10'd27, 10'd17};
parameter Y27X18={10'd27, 10'd18};
parameter Y27X19={10'd27, 10'd19};
parameter Y27X20={10'd27, 10'd20};
parameter Y27X21={10'd27, 10'd21};
parameter Y27X22={10'd27, 10'd22};
parameter Y27X23={10'd27, 10'd23};
parameter Y27X24={10'd27, 10'd24};
parameter Y27X25={10'd27, 10'd25};
parameter Y27X26={10'd27, 10'd26};
parameter Y27X27={10'd27, 10'd27};
parameter Y27X28={10'd27, 10'd28};
parameter Y28X1={10'd28, 10'd1};
parameter Y28X2={10'd28, 10'd2};
parameter Y28X3={10'd28, 10'd3};
parameter Y28X4={10'd28, 10'd4};
parameter Y28X5={10'd28, 10'd5};
parameter Y28X6={10'd28, 10'd6};
parameter Y28X7={10'd28, 10'd7};
parameter Y28X8={10'd28, 10'd8};
parameter Y28X9={10'd28, 10'd9};
parameter Y28X10={10'd28, 10'd10};
parameter Y28X11={10'd28, 10'd11};
parameter Y28X12={10'd28, 10'd12};
parameter Y28X13={10'd28, 10'd13};
parameter Y28X14={10'd28, 10'd14};
parameter Y28X15={10'd28, 10'd15};
parameter Y28X16={10'd28, 10'd16};
parameter Y28X17={10'd28, 10'd17};
parameter Y28X18={10'd28, 10'd18};
parameter Y28X19={10'd28, 10'd19};
parameter Y28X20={10'd28, 10'd20};
parameter Y28X21={10'd28, 10'd21};
parameter Y28X22={10'd28, 10'd22};
parameter Y28X23={10'd28, 10'd23};
parameter Y28X24={10'd28, 10'd24};
parameter Y28X25={10'd28, 10'd25};
parameter Y28X26={10'd28, 10'd26};
parameter Y28X27={10'd28, 10'd27};
parameter Y28X28={10'd28, 10'd28};
parameter Y29X1={10'd29, 10'd1};
parameter Y29X2={10'd29, 10'd2};
parameter Y29X3={10'd29, 10'd3};
parameter Y29X4={10'd29, 10'd4};
parameter Y29X5={10'd29, 10'd5};
parameter Y29X6={10'd29, 10'd6};
parameter Y29X7={10'd29, 10'd7};
parameter Y29X8={10'd29, 10'd8};
parameter Y29X9={10'd29, 10'd9};
parameter Y29X10={10'd29, 10'd10};
parameter Y29X11={10'd29, 10'd11};
parameter Y29X12={10'd29, 10'd12};
parameter Y29X13={10'd29, 10'd13};
parameter Y29X14={10'd29, 10'd14};
parameter Y29X15={10'd29, 10'd15};
parameter Y29X16={10'd29, 10'd16};
parameter Y29X17={10'd29, 10'd17};
parameter Y29X18={10'd29, 10'd18};
parameter Y29X19={10'd29, 10'd19};
parameter Y29X20={10'd29, 10'd20};
parameter Y29X21={10'd29, 10'd21};
parameter Y29X22={10'd29, 10'd22};
parameter Y29X23={10'd29, 10'd23};
parameter Y29X24={10'd29, 10'd24};
parameter Y29X25={10'd29, 10'd25};
parameter Y29X26={10'd29, 10'd26};
parameter Y29X27={10'd29, 10'd27};
parameter Y29X28={10'd29, 10'd28};
parameter Y30X1={10'd30, 10'd1};
parameter Y30X2={10'd30, 10'd2};
parameter Y30X3={10'd30, 10'd3};
parameter Y30X4={10'd30, 10'd4};
parameter Y30X5={10'd30, 10'd5};
parameter Y30X6={10'd30, 10'd6};
parameter Y30X7={10'd30, 10'd7};
parameter Y30X8={10'd30, 10'd8};
parameter Y30X9={10'd30, 10'd9};
parameter Y30X10={10'd30, 10'd10};
parameter Y30X11={10'd30, 10'd11};
parameter Y30X12={10'd30, 10'd12};
parameter Y30X13={10'd30, 10'd13};
parameter Y30X14={10'd30, 10'd14};
parameter Y30X15={10'd30, 10'd15};
parameter Y30X16={10'd30, 10'd16};
parameter Y30X17={10'd30, 10'd17};
parameter Y30X18={10'd30, 10'd18};
parameter Y30X19={10'd30, 10'd19};
parameter Y30X20={10'd30, 10'd20};
parameter Y30X21={10'd30, 10'd21};
parameter Y30X22={10'd30, 10'd22};
parameter Y30X23={10'd30, 10'd23};
parameter Y30X24={10'd30, 10'd24};
parameter Y30X25={10'd30, 10'd25};
parameter Y30X26={10'd30, 10'd26};
parameter Y30X27={10'd30, 10'd27};
parameter Y30X28={10'd30, 10'd28};
parameter Y31X1={10'd31, 10'd1};
parameter Y31X2={10'd31, 10'd2};
parameter Y31X3={10'd31, 10'd3};
parameter Y31X4={10'd31, 10'd4};
parameter Y31X5={10'd31, 10'd5};
parameter Y31X6={10'd31, 10'd6};
parameter Y31X7={10'd31, 10'd7};
parameter Y31X8={10'd31, 10'd8};
parameter Y31X9={10'd31, 10'd9};
parameter Y31X10={10'd31, 10'd10};
parameter Y31X11={10'd31, 10'd11};
parameter Y31X12={10'd31, 10'd12};
parameter Y31X13={10'd31, 10'd13};
parameter Y31X14={10'd31, 10'd14};
parameter Y31X15={10'd31, 10'd15};
parameter Y31X16={10'd31, 10'd16};
parameter Y31X17={10'd31, 10'd17};
parameter Y31X18={10'd31, 10'd18};
parameter Y31X19={10'd31, 10'd19};
parameter Y31X20={10'd31, 10'd20};
parameter Y31X21={10'd31, 10'd21};
parameter Y31X22={10'd31, 10'd22};
parameter Y31X23={10'd31, 10'd23};
parameter Y31X24={10'd31, 10'd24};
parameter Y31X25={10'd31, 10'd25};
parameter Y31X26={10'd31, 10'd26};
parameter Y31X27={10'd31, 10'd27};
parameter Y31X28={10'd31, 10'd28};
parameter Y32X1={10'd32, 10'd1};
parameter Y32X2={10'd32, 10'd2};
parameter Y32X3={10'd32, 10'd3};
parameter Y32X4={10'd32, 10'd4};
parameter Y32X5={10'd32, 10'd5};
parameter Y32X6={10'd32, 10'd6};
parameter Y32X7={10'd32, 10'd7};
parameter Y32X8={10'd32, 10'd8};
parameter Y32X9={10'd32, 10'd9};
parameter Y32X10={10'd32, 10'd10};
parameter Y32X11={10'd32, 10'd11};
parameter Y32X12={10'd32, 10'd12};
parameter Y32X13={10'd32, 10'd13};
parameter Y32X14={10'd32, 10'd14};
parameter Y32X15={10'd32, 10'd15};
parameter Y32X16={10'd32, 10'd16};
parameter Y32X17={10'd32, 10'd17};
parameter Y32X18={10'd32, 10'd18};
parameter Y32X19={10'd32, 10'd19};
parameter Y32X20={10'd32, 10'd20};
parameter Y32X21={10'd32, 10'd21};
parameter Y32X22={10'd32, 10'd22};
parameter Y32X23={10'd32, 10'd23};
parameter Y32X24={10'd32, 10'd24};
parameter Y32X25={10'd32, 10'd25};
parameter Y32X26={10'd32, 10'd26};
parameter Y32X27={10'd32, 10'd27};
parameter Y32X28={10'd32, 10'd28};
parameter Y33X1={10'd33, 10'd1};
parameter Y33X2={10'd33, 10'd2};
parameter Y33X3={10'd33, 10'd3};
parameter Y33X4={10'd33, 10'd4};
parameter Y33X5={10'd33, 10'd5};
parameter Y33X6={10'd33, 10'd6};
parameter Y33X7={10'd33, 10'd7};
parameter Y33X8={10'd33, 10'd8};
parameter Y33X9={10'd33, 10'd9};
parameter Y33X10={10'd33, 10'd10};
parameter Y33X11={10'd33, 10'd11};
parameter Y33X12={10'd33, 10'd12};
parameter Y33X13={10'd33, 10'd13};
parameter Y33X14={10'd33, 10'd14};
parameter Y33X15={10'd33, 10'd15};
parameter Y33X16={10'd33, 10'd16};
parameter Y33X17={10'd33, 10'd17};
parameter Y33X18={10'd33, 10'd18};
parameter Y33X19={10'd33, 10'd19};
parameter Y33X20={10'd33, 10'd20};
parameter Y33X21={10'd33, 10'd21};
parameter Y33X22={10'd33, 10'd22};
parameter Y33X23={10'd33, 10'd23};
parameter Y33X24={10'd33, 10'd24};
parameter Y33X25={10'd33, 10'd25};
parameter Y33X26={10'd33, 10'd26};
parameter Y33X27={10'd33, 10'd27};
parameter Y33X28={10'd33, 10'd28};
parameter Y34X1={10'd34, 10'd1};
parameter Y34X2={10'd34, 10'd2};
parameter Y34X3={10'd34, 10'd3};
parameter Y34X4={10'd34, 10'd4};
parameter Y34X5={10'd34, 10'd5};
parameter Y34X6={10'd34, 10'd6};
parameter Y34X7={10'd34, 10'd7};
parameter Y34X8={10'd34, 10'd8};
parameter Y34X9={10'd34, 10'd9};
parameter Y34X10={10'd34, 10'd10};
parameter Y34X11={10'd34, 10'd11};
parameter Y34X12={10'd34, 10'd12};
parameter Y34X13={10'd34, 10'd13};
parameter Y34X14={10'd34, 10'd14};
parameter Y34X15={10'd34, 10'd15};
parameter Y34X16={10'd34, 10'd16};
parameter Y34X17={10'd34, 10'd17};
parameter Y34X18={10'd34, 10'd18};
parameter Y34X19={10'd34, 10'd19};
parameter Y34X20={10'd34, 10'd20};
parameter Y34X21={10'd34, 10'd21};
parameter Y34X22={10'd34, 10'd22};
parameter Y34X23={10'd34, 10'd23};
parameter Y34X24={10'd34, 10'd24};
parameter Y34X25={10'd34, 10'd25};
parameter Y34X26={10'd34, 10'd26};
parameter Y34X27={10'd34, 10'd27};
parameter Y34X28={10'd34, 10'd28};
parameter Y35X1={10'd35, 10'd1};
parameter Y35X2={10'd35, 10'd2};
parameter Y35X3={10'd35, 10'd3};
parameter Y35X4={10'd35, 10'd4};
parameter Y35X5={10'd35, 10'd5};
parameter Y35X6={10'd35, 10'd6};
parameter Y35X7={10'd35, 10'd7};
parameter Y35X8={10'd35, 10'd8};
parameter Y35X9={10'd35, 10'd9};
parameter Y35X10={10'd35, 10'd10};
parameter Y35X11={10'd35, 10'd11};
parameter Y35X12={10'd35, 10'd12};
parameter Y35X13={10'd35, 10'd13};
parameter Y35X14={10'd35, 10'd14};
parameter Y35X15={10'd35, 10'd15};
parameter Y35X16={10'd35, 10'd16};
parameter Y35X17={10'd35, 10'd17};
parameter Y35X18={10'd35, 10'd18};
parameter Y35X19={10'd35, 10'd19};
parameter Y35X20={10'd35, 10'd20};
parameter Y35X21={10'd35, 10'd21};
parameter Y35X22={10'd35, 10'd22};
parameter Y35X23={10'd35, 10'd23};
parameter Y35X24={10'd35, 10'd24};
parameter Y35X25={10'd35, 10'd25};
parameter Y35X26={10'd35, 10'd26};
parameter Y35X27={10'd35, 10'd27};
parameter Y35X28={10'd35, 10'd28};

parameter YY0XX0={4'd15,4'd0,4'd0};
parameter YY0XX1={4'd3,4'd3,4'd3};
parameter YY0XX2={4'd6,4'd5,4'd5};
parameter YY0XX3={4'd6,4'd6,4'd5};
parameter YY0XX4={4'd7,4'd7,4'd6};
parameter YY0XX5={4'd15,4'd0,4'd0};
parameter YY0XX6={4'd15,4'd0,4'd0};
parameter YY0XX7={4'd15,4'd0,4'd0};
parameter YY0XX8={4'd15,4'd0,4'd0};
parameter YY0XX9={4'd15,4'd0,4'd0};
parameter YY0XX10={4'd15,4'd0,4'd0};
parameter YY0XX11={4'd15,4'd0,4'd0};
parameter YY0XX12={4'd15,4'd0,4'd0};
parameter YY0XX13={4'd15,4'd0,4'd0};
parameter YY0XX14={4'd15,4'd0,4'd0};
parameter YY0XX15={4'd15,4'd0,4'd0};
parameter YY0XX16={4'd15,4'd0,4'd0};
parameter YY0XX17={4'd15,4'd0,4'd0};
parameter YY0XX18={4'd15,4'd0,4'd0};
parameter YY0XX19={4'd15,4'd0,4'd0};
parameter YY0XX20={4'd15,4'd0,4'd0};
parameter YY0XX21={4'd15,4'd0,4'd0};
parameter YY0XX22={4'd15,4'd0,4'd0};
parameter YY0XX23={4'd15,4'd0,4'd0};
parameter YY0XX24={4'd15,4'd0,4'd0};
parameter YY0XX25={4'd15,4'd0,4'd0};
parameter YY0XX26={4'd15,4'd0,4'd0};
parameter YY0XX27={4'd15,4'd0,4'd0};
parameter YY0XX28={4'd15,4'd0,4'd0};
parameter YY1XX1={4'd8,4'd8,4'd8};
parameter YY1XX2={4'd12,4'd12,4'd12};
parameter YY1XX3={4'd13,4'd12,4'd12};
parameter YY1XX4={4'd13,4'd13,4'd13};
parameter YY1XX5={4'd11,4'd11,4'd10};
parameter YY1XX6={4'd8,4'd8,4'd7};
parameter YY1XX7={4'd15,4'd0,4'd0};
parameter YY1XX8={4'd15,4'd0,4'd0};
parameter YY1XX9={4'd15,4'd0,4'd0};
parameter YY1XX10={4'd15,4'd0,4'd0};
parameter YY1XX11={4'd15,4'd0,4'd0};
parameter YY1XX12={4'd15,4'd0,4'd0};
parameter YY1XX13={4'd15,4'd0,4'd0};
parameter YY1XX14={4'd15,4'd0,4'd0};
parameter YY1XX15={4'd15,4'd0,4'd0};
parameter YY1XX16={4'd15,4'd0,4'd0};
parameter YY1XX17={4'd15,4'd0,4'd0};
parameter YY1XX18={4'd15,4'd0,4'd0};
parameter YY1XX19={4'd15,4'd0,4'd0};
parameter YY1XX20={4'd15,4'd0,4'd0};
parameter YY1XX21={4'd15,4'd0,4'd0};
parameter YY1XX22={4'd15,4'd0,4'd0};
parameter YY1XX23={4'd15,4'd0,4'd0};
parameter YY1XX24={4'd15,4'd0,4'd0};
parameter YY1XX25={4'd15,4'd0,4'd0};
parameter YY1XX26={4'd15,4'd0,4'd0};
parameter YY1XX27={4'd15,4'd0,4'd0};
parameter YY1XX28={4'd15,4'd0,4'd0};
parameter YY2XX1={4'd11,4'd11,4'd11};
parameter YY2XX2={4'd15,4'd15,4'd15};
parameter YY2XX3={4'd15,4'd15,4'd15};
parameter YY2XX4={4'd15,4'd15,4'd15};
parameter YY2XX5={4'd15,4'd15,4'd15};
parameter YY2XX6={4'd14,4'd13,4'd13};
parameter YY2XX7={4'd10,4'd9,4'd9};
parameter YY2XX8={4'd15,4'd0,4'd0};
parameter YY2XX9={4'd15,4'd0,4'd0};
parameter YY2XX10={4'd15,4'd0,4'd0};
parameter YY2XX11={4'd15,4'd0,4'd0};
parameter YY2XX12={4'd15,4'd0,4'd0};
parameter YY2XX13={4'd15,4'd0,4'd0};
parameter YY2XX14={4'd15,4'd0,4'd0};
parameter YY2XX15={4'd15,4'd0,4'd0};
parameter YY2XX16={4'd15,4'd0,4'd0};
parameter YY2XX17={4'd15,4'd0,4'd0};
parameter YY2XX18={4'd15,4'd0,4'd0};
parameter YY2XX19={4'd15,4'd0,4'd0};
parameter YY2XX20={4'd15,4'd0,4'd0};
parameter YY2XX21={4'd15,4'd0,4'd0};
parameter YY2XX22={4'd15,4'd0,4'd0};
parameter YY2XX23={4'd15,4'd0,4'd0};
parameter YY2XX24={4'd15,4'd0,4'd0};
parameter YY2XX25={4'd15,4'd0,4'd0};
parameter YY2XX26={4'd15,4'd0,4'd0};
parameter YY2XX27={4'd15,4'd0,4'd0};
parameter YY2XX28={4'd15,4'd0,4'd0};
parameter YY3XX1={4'd11,4'd11,4'd11};
parameter YY3XX2={4'd15,4'd15,4'd15};
parameter YY3XX3={4'd15,4'd15,4'd15};
parameter YY3XX4={4'd15,4'd15,4'd15};
parameter YY3XX5={4'd15,4'd15,4'd15};
parameter YY3XX6={4'd15,4'd15,4'd15};
parameter YY3XX7={4'd15,4'd14,4'd15};
parameter YY3XX8={4'd12,4'd11,4'd11};
parameter YY3XX9={4'd15,4'd0,4'd0};
parameter YY3XX10={4'd15,4'd0,4'd0};
parameter YY3XX11={4'd15,4'd0,4'd0};
parameter YY3XX12={4'd15,4'd0,4'd0};
parameter YY3XX13={4'd15,4'd0,4'd0};
parameter YY3XX14={4'd15,4'd0,4'd0};
parameter YY3XX15={4'd15,4'd0,4'd0};
parameter YY3XX16={4'd15,4'd0,4'd0};
parameter YY3XX17={4'd15,4'd0,4'd0};
parameter YY3XX18={4'd15,4'd0,4'd0};
parameter YY3XX19={4'd15,4'd0,4'd0};
parameter YY3XX20={4'd15,4'd0,4'd0};
parameter YY3XX21={4'd15,4'd0,4'd0};
parameter YY3XX22={4'd15,4'd0,4'd0};
parameter YY3XX23={4'd15,4'd0,4'd0};
parameter YY3XX24={4'd15,4'd0,4'd0};
parameter YY3XX25={4'd15,4'd0,4'd0};
parameter YY3XX26={4'd15,4'd0,4'd0};
parameter YY3XX27={4'd15,4'd0,4'd0};
parameter YY3XX28={4'd15,4'd0,4'd0};
parameter YY4XX1={4'd10,4'd10,4'd10};
parameter YY4XX2={4'd13,4'd13,4'd14};
parameter YY4XX3={4'd15,4'd15,4'd15};
parameter YY4XX4={4'd15,4'd15,4'd15};
parameter YY4XX5={4'd15,4'd15,4'd15};
parameter YY4XX6={4'd15,4'd15,4'd15};
parameter YY4XX7={4'd15,4'd15,4'd15};
parameter YY4XX8={4'd15,4'd15,4'd15};
parameter YY4XX9={4'd13,4'd12,4'd11};
parameter YY4XX10={4'd15,4'd0,4'd0};
parameter YY4XX11={4'd15,4'd0,4'd0};
parameter YY4XX12={4'd15,4'd0,4'd0};
parameter YY4XX13={4'd15,4'd0,4'd0};
parameter YY4XX14={4'd15,4'd0,4'd0};
parameter YY4XX15={4'd15,4'd0,4'd0};
parameter YY4XX16={4'd15,4'd0,4'd0};
parameter YY4XX17={4'd15,4'd0,4'd0};
parameter YY4XX18={4'd15,4'd0,4'd0};
parameter YY4XX19={4'd15,4'd0,4'd0};
parameter YY4XX20={4'd15,4'd0,4'd0};
parameter YY4XX21={4'd15,4'd0,4'd0};
parameter YY4XX22={4'd15,4'd0,4'd0};
parameter YY4XX23={4'd15,4'd0,4'd0};
parameter YY4XX24={4'd15,4'd0,4'd0};
parameter YY4XX25={4'd15,4'd0,4'd0};
parameter YY4XX26={4'd15,4'd0,4'd0};
parameter YY4XX27={4'd15,4'd0,4'd0};
parameter YY4XX28={4'd15,4'd0,4'd0};
parameter YY5XX1={4'd7,4'd8,4'd7};
parameter YY5XX2={4'd11,4'd11,4'd11};
parameter YY5XX3={4'd14,4'd14,4'd14};
parameter YY5XX4={4'd15,4'd15,4'd15};
parameter YY5XX5={4'd15,4'd15,4'd15};
parameter YY5XX6={4'd15,4'd15,4'd15};
parameter YY5XX7={4'd15,4'd15,4'd15};
parameter YY5XX8={4'd15,4'd15,4'd15};
parameter YY5XX9={4'd15,4'd15,4'd15};
parameter YY5XX10={4'd13,4'd12,4'd12};
parameter YY5XX11={4'd15,4'd0,4'd0};
parameter YY5XX12={4'd15,4'd0,4'd0};
parameter YY5XX13={4'd15,4'd0,4'd0};
parameter YY5XX14={4'd15,4'd0,4'd0};
parameter YY5XX15={4'd15,4'd0,4'd0};
parameter YY5XX16={4'd15,4'd0,4'd0};
parameter YY5XX17={4'd15,4'd0,4'd0};
parameter YY5XX18={4'd15,4'd0,4'd0};
parameter YY5XX19={4'd15,4'd0,4'd0};
parameter YY5XX20={4'd15,4'd0,4'd0};
parameter YY5XX21={4'd15,4'd0,4'd0};
parameter YY5XX22={4'd15,4'd0,4'd0};
parameter YY5XX23={4'd15,4'd0,4'd0};
parameter YY5XX24={4'd15,4'd0,4'd0};
parameter YY5XX25={4'd15,4'd0,4'd0};
parameter YY5XX26={4'd15,4'd0,4'd0};
parameter YY5XX27={4'd15,4'd0,4'd0};
parameter YY5XX28={4'd15,4'd0,4'd0};
parameter YY6XX1={4'd5,4'd5,4'd5};
parameter YY6XX2={4'd8,4'd9,4'd9};
parameter YY6XX3={4'd12,4'd12,4'd12};
parameter YY6XX4={4'd15,4'd15,4'd15};
parameter YY6XX5={4'd15,4'd15,4'd15};
parameter YY6XX6={4'd15,4'd15,4'd15};
parameter YY6XX7={4'd15,4'd15,4'd15};
parameter YY6XX8={4'd15,4'd15,4'd15};
parameter YY6XX9={4'd15,4'd15,4'd15};
parameter YY6XX10={4'd15,4'd14,4'd15};
parameter YY6XX11={4'd13,4'd12,4'd13};
parameter YY6XX12={4'd10,4'd10,4'd10};
parameter YY6XX13={4'd15,4'd0,4'd0};
parameter YY6XX14={4'd15,4'd0,4'd0};
parameter YY6XX15={4'd15,4'd0,4'd0};
parameter YY6XX16={4'd15,4'd0,4'd0};
parameter YY6XX17={4'd15,4'd0,4'd0};
parameter YY6XX18={4'd15,4'd0,4'd0};
parameter YY6XX19={4'd4,4'd3,4'd3};
parameter YY6XX20={4'd4,4'd3,4'd3};
parameter YY6XX21={4'd3,4'd3,4'd2};
parameter YY6XX22={4'd15,4'd0,4'd0};
parameter YY6XX23={4'd15,4'd0,4'd0};
parameter YY6XX24={4'd15,4'd0,4'd0};
parameter YY6XX25={4'd15,4'd0,4'd0};
parameter YY6XX26={4'd15,4'd0,4'd0};
parameter YY6XX27={4'd15,4'd0,4'd0};
parameter YY6XX28={4'd15,4'd0,4'd0};
parameter YY7XX1={4'd15,4'd0,4'd0};
parameter YY7XX2={4'd5,4'd5,4'd5};
parameter YY7XX3={4'd8,4'd8,4'd9};
parameter YY7XX4={4'd12,4'd12,4'd12};
parameter YY7XX5={4'd14,4'd14,4'd14};
parameter YY7XX6={4'd15,4'd15,4'd15};
parameter YY7XX7={4'd15,4'd15,4'd15};
parameter YY7XX8={4'd15,4'd15,4'd15};
parameter YY7XX9={4'd15,4'd15,4'd15};
parameter YY7XX10={4'd15,4'd15,4'd15};
parameter YY7XX11={4'd15,4'd15,4'd15};
parameter YY7XX12={4'd15,4'd14,4'd14};
parameter YY7XX13={4'd11,4'd11,4'd11};
parameter YY7XX14={4'd15,4'd0,4'd0};
parameter YY7XX15={4'd15,4'd0,4'd0};
parameter YY7XX16={4'd15,4'd0,4'd0};
parameter YY7XX17={4'd15,4'd0,4'd0};
parameter YY7XX18={4'd7,4'd6,4'd6};
parameter YY7XX19={4'd9,4'd9,4'd8};
parameter YY7XX20={4'd10,4'd9,4'd9};
parameter YY7XX21={4'd7,4'd7,4'd7};
parameter YY7XX22={4'd4,4'd4,4'd3};
parameter YY7XX23={4'd15,4'd0,4'd0};
parameter YY7XX24={4'd15,4'd0,4'd0};
parameter YY7XX25={4'd15,4'd0,4'd0};
parameter YY7XX26={4'd15,4'd0,4'd0};
parameter YY7XX27={4'd15,4'd0,4'd0};
parameter YY7XX28={4'd15,4'd0,4'd0};
parameter YY8XX1={4'd15,4'd0,4'd0};
parameter YY8XX2={4'd15,4'd0,4'd0};
parameter YY8XX3={4'd4,4'd4,4'd4};
parameter YY8XX4={4'd8,4'd7,4'd8};
parameter YY8XX5={4'd11,4'd10,4'd11};
parameter YY8XX6={4'd14,4'd14,4'd14};
parameter YY8XX7={4'd15,4'd15,4'd15};
parameter YY8XX8={4'd15,4'd15,4'd15};
parameter YY8XX9={4'd15,4'd15,4'd15};
parameter YY8XX10={4'd15,4'd15,4'd15};
parameter YY8XX11={4'd15,4'd15,4'd15};
parameter YY8XX12={4'd15,4'd15,4'd15};
parameter YY8XX13={4'd14,4'd14,4'd14};
parameter YY8XX14={4'd12,4'd11,4'd11};
parameter YY8XX15={4'd9,4'd8,4'd8};
parameter YY8XX16={4'd7,4'd7,4'd7};
parameter YY8XX17={4'd7,4'd6,4'd6};
parameter YY8XX18={4'd9,4'd8,4'd8};
parameter YY8XX19={4'd13,4'd12,4'd12};
parameter YY8XX20={4'd15,4'd14,4'd14};
parameter YY8XX21={4'd12,4'd12,4'd11};
parameter YY8XX22={4'd8,4'd7,4'd7};
parameter YY8XX23={4'd9,4'd8,4'd7};
parameter YY8XX24={4'd15,4'd0,4'd0};
parameter YY8XX25={4'd15,4'd0,4'd0};
parameter YY8XX26={4'd15,4'd0,4'd0};
parameter YY8XX27={4'd15,4'd0,4'd0};
parameter YY8XX28={4'd15,4'd0,4'd0};
parameter YY9XX1={4'd15,4'd0,4'd0};
parameter YY9XX2={4'd15,4'd0,4'd0};
parameter YY9XX3={4'd15,4'd0,4'd0};
parameter YY9XX4={4'd4,4'd3,4'd4};
parameter YY9XX5={4'd7,4'd6,4'd7};
parameter YY9XX6={4'd11,4'd10,4'd11};
parameter YY9XX7={4'd14,4'd14,4'd14};
parameter YY9XX8={4'd15,4'd15,4'd15};
parameter YY9XX9={4'd15,4'd15,4'd15};
parameter YY9XX10={4'd15,4'd15,4'd15};
parameter YY9XX11={4'd15,4'd15,4'd15};
parameter YY9XX12={4'd15,4'd15,4'd15};
parameter YY9XX13={4'd15,4'd15,4'd15};
parameter YY9XX14={4'd15,4'd15,4'd15};
parameter YY9XX15={4'd13,4'd13,4'd13};
parameter YY9XX16={4'd12,4'd11,4'd11};
parameter YY9XX17={4'd10,4'd10,4'd10};
parameter YY9XX18={4'd11,4'd10,4'd10};
parameter YY9XX19={4'd14,4'd13,4'd13};
parameter YY9XX20={4'd15,4'd15,4'd15};
parameter YY9XX21={4'd15,4'd14,4'd14};
parameter YY9XX22={4'd12,4'd12,4'd11};
parameter YY9XX23={4'd9,4'd8,4'd7};
parameter YY9XX24={4'd8,4'd7,4'd6};
parameter YY9XX25={4'd15,4'd0,4'd0};
parameter YY9XX26={4'd15,4'd0,4'd0};
parameter YY9XX27={4'd15,4'd0,4'd0};
parameter YY9XX28={4'd15,4'd0,4'd0};
parameter YY10XX1={4'd15,4'd0,4'd0};
parameter YY10XX2={4'd15,4'd0,4'd0};
parameter YY10XX3={4'd15,4'd0,4'd0};
parameter YY10XX4={4'd15,4'd0,4'd0};
parameter YY10XX5={4'd5,4'd4,4'd5};
parameter YY10XX6={4'd8,4'd7,4'd8};
parameter YY10XX7={4'd11,4'd11,4'd11};
parameter YY10XX8={4'd13,4'd13,4'd13};
parameter YY10XX9={4'd15,4'd15,4'd15};
parameter YY10XX10={4'd15,4'd15,4'd15};
parameter YY10XX11={4'd15,4'd15,4'd15};
parameter YY10XX12={4'd15,4'd15,4'd15};
parameter YY10XX13={4'd15,4'd15,4'd15};
parameter YY10XX14={4'd15,4'd15,4'd15};
parameter YY10XX15={4'd15,4'd15,4'd15};
parameter YY10XX16={4'd15,4'd15,4'd15};
parameter YY10XX17={4'd14,4'd14,4'd14};
parameter YY10XX18={4'd13,4'd13,4'd13};
parameter YY10XX19={4'd14,4'd13,4'd13};
parameter YY10XX20={4'd15,4'd15,4'd15};
parameter YY10XX21={4'd15,4'd15,4'd15};
parameter YY10XX22={4'd15,4'd15,4'd15};
parameter YY10XX23={4'd12,4'd11,4'd10};
parameter YY10XX24={4'd9,4'd8,4'd7};
parameter YY10XX25={4'd15,4'd0,4'd0};
parameter YY10XX26={4'd15,4'd0,4'd0};
parameter YY10XX27={4'd15,4'd0,4'd0};
parameter YY10XX28={4'd15,4'd0,4'd0};
parameter YY11XX1={4'd15,4'd0,4'd0};
parameter YY11XX2={4'd15,4'd0,4'd0};
parameter YY11XX3={4'd15,4'd0,4'd0};
parameter YY11XX4={4'd4,4'd3,4'd4};
parameter YY11XX5={4'd6,4'd5,4'd6};
parameter YY11XX6={4'd9,4'd9,4'd9};
parameter YY11XX7={4'd12,4'd11,4'd12};
parameter YY11XX8={4'd13,4'd13,4'd13};
parameter YY11XX9={4'd15,4'd15,4'd15};
parameter YY11XX10={4'd15,4'd15,4'd15};
parameter YY11XX11={4'd15,4'd15,4'd15};
parameter YY11XX12={4'd15,4'd15,4'd15};
parameter YY11XX13={4'd15,4'd15,4'd15};
parameter YY11XX14={4'd15,4'd15,4'd15};
parameter YY11XX15={4'd15,4'd15,4'd15};
parameter YY11XX16={4'd15,4'd15,4'd15};
parameter YY11XX17={4'd15,4'd15,4'd15};
parameter YY11XX18={4'd14,4'd14,4'd14};
parameter YY11XX19={4'd14,4'd13,4'd14};
parameter YY11XX20={4'd14,4'd14,4'd14};
parameter YY11XX21={4'd15,4'd15,4'd15};
parameter YY11XX22={4'd15,4'd15,4'd15};
parameter YY11XX23={4'd15,4'd15,4'd14};
parameter YY11XX24={4'd13,4'd12,4'd11};
parameter YY11XX25={4'd7,4'd6,4'd5};
parameter YY11XX26={4'd15,4'd0,4'd0};
parameter YY11XX27={4'd15,4'd0,4'd0};
parameter YY11XX28={4'd15,4'd0,4'd0};
parameter YY12XX1={4'd15,4'd0,4'd0};
parameter YY12XX2={4'd15,4'd0,4'd0};
parameter YY12XX3={4'd3,4'd2,4'd3};
parameter YY12XX4={4'd5,4'd5,4'd5};
parameter YY12XX5={4'd8,4'd8,4'd8};
parameter YY12XX6={4'd12,4'd12,4'd12};
parameter YY12XX7={4'd15,4'd14,4'd15};
parameter YY12XX8={4'd15,4'd14,4'd15};
parameter YY12XX9={4'd15,4'd15,4'd15};
parameter YY12XX10={4'd15,4'd15,4'd15};
parameter YY12XX11={4'd15,4'd15,4'd15};
parameter YY12XX12={4'd15,4'd15,4'd15};
parameter YY12XX13={4'd15,4'd15,4'd15};
parameter YY12XX14={4'd15,4'd15,4'd15};
parameter YY12XX15={4'd15,4'd15,4'd15};
parameter YY12XX16={4'd15,4'd15,4'd15};
parameter YY12XX17={4'd15,4'd15,4'd15};
parameter YY12XX18={4'd15,4'd15,4'd15};
parameter YY12XX19={4'd15,4'd15,4'd15};
parameter YY12XX20={4'd15,4'd15,4'd15};
parameter YY12XX21={4'd15,4'd15,4'd15};
parameter YY12XX22={4'd15,4'd15,4'd15};
parameter YY12XX23={4'd15,4'd15,4'd15};
parameter YY12XX24={4'd15,4'd15,4'd14};
parameter YY12XX25={4'd10,4'd10,4'd9};
parameter YY12XX26={4'd15,4'd0,4'd0};
parameter YY12XX27={4'd15,4'd0,4'd0};
parameter YY12XX28={4'd15,4'd0,4'd0};
parameter YY13XX1={4'd15,4'd0,4'd0};
parameter YY13XX2={4'd15,4'd0,4'd0};
parameter YY13XX3={4'd6,4'd6,4'd6};
parameter YY13XX4={4'd9,4'd9,4'd9};
parameter YY13XX5={4'd12,4'd12,4'd12};
parameter YY13XX6={4'd14,4'd14,4'd14};
parameter YY13XX7={4'd15,4'd15,4'd15};
parameter YY13XX8={4'd15,4'd15,4'd15};
parameter YY13XX9={4'd15,4'd15,4'd15};
parameter YY13XX10={4'd15,4'd15,4'd15};
parameter YY13XX11={4'd15,4'd15,4'd15};
parameter YY13XX12={4'd15,4'd15,4'd15};
parameter YY13XX13={4'd15,4'd15,4'd15};
parameter YY13XX14={4'd15,4'd15,4'd15};
parameter YY13XX15={4'd15,4'd15,4'd15};
parameter YY13XX16={4'd15,4'd15,4'd15};
parameter YY13XX17={4'd15,4'd15,4'd15};
parameter YY13XX18={4'd15,4'd15,4'd15};
parameter YY13XX19={4'd15,4'd15,4'd15};
parameter YY13XX20={4'd15,4'd15,4'd15};
parameter YY13XX21={4'd15,4'd15,4'd15};
parameter YY13XX22={4'd15,4'd15,4'd15};
parameter YY13XX23={4'd15,4'd15,4'd15};
parameter YY13XX24={4'd15,4'd14,4'd14};
parameter YY13XX25={4'd11,4'd10,4'd9};
parameter YY13XX26={4'd15,4'd0,4'd0};
parameter YY13XX27={4'd15,4'd0,4'd0};
parameter YY13XX28={4'd15,4'd0,4'd0};
parameter YY14XX1={4'd15,4'd0,4'd0};
parameter YY14XX2={4'd5,4'd5,4'd5};
parameter YY14XX3={4'd8,4'd8,4'd8};
parameter YY14XX4={4'd12,4'd12,4'd12};
parameter YY14XX5={4'd14,4'd14,4'd14};
parameter YY14XX6={4'd15,4'd15,4'd15};
parameter YY14XX7={4'd15,4'd15,4'd15};
parameter YY14XX8={4'd15,4'd15,4'd15};
parameter YY14XX9={4'd15,4'd15,4'd15};
parameter YY14XX10={4'd15,4'd15,4'd15};
parameter YY14XX11={4'd15,4'd15,4'd15};
parameter YY14XX12={4'd15,4'd15,4'd15};
parameter YY14XX13={4'd15,4'd15,4'd15};
parameter YY14XX14={4'd15,4'd15,4'd15};
parameter YY14XX15={4'd15,4'd15,4'd15};
parameter YY14XX16={4'd15,4'd15,4'd15};
parameter YY14XX17={4'd15,4'd15,4'd15};
parameter YY14XX18={4'd15,4'd15,4'd15};
parameter YY14XX19={4'd15,4'd15,4'd15};
parameter YY14XX20={4'd15,4'd15,4'd15};
parameter YY14XX21={4'd15,4'd15,4'd15};
parameter YY14XX22={4'd15,4'd15,4'd15};
parameter YY14XX23={4'd15,4'd15,4'd15};
parameter YY14XX24={4'd15,4'd15,4'd14};
parameter YY14XX25={4'd11,4'd10,4'd10};
parameter YY14XX26={4'd15,4'd0,4'd0};
parameter YY14XX27={4'd15,4'd0,4'd0};
parameter YY14XX28={4'd15,4'd0,4'd0};
parameter YY15XX1={4'd15,4'd0,4'd0};
parameter YY15XX2={4'd6,4'd6,4'd5};
parameter YY15XX3={4'd9,4'd10,4'd9};
parameter YY15XX4={4'd13,4'd14,4'd13};
parameter YY15XX5={4'd15,4'd15,4'd15};
parameter YY15XX6={4'd15,4'd15,4'd15};
parameter YY15XX7={4'd15,4'd15,4'd15};
parameter YY15XX8={4'd15,4'd15,4'd15};
parameter YY15XX9={4'd15,4'd15,4'd15};
parameter YY15XX10={4'd15,4'd15,4'd15};
parameter YY15XX11={4'd15,4'd15,4'd15};
parameter YY15XX12={4'd15,4'd15,4'd15};
parameter YY15XX13={4'd15,4'd15,4'd15};
parameter YY15XX14={4'd15,4'd15,4'd15};
parameter YY15XX15={4'd15,4'd15,4'd15};
parameter YY15XX16={4'd15,4'd15,4'd15};
parameter YY15XX17={4'd15,4'd15,4'd15};
parameter YY15XX18={4'd15,4'd15,4'd15};
parameter YY15XX19={4'd15,4'd15,4'd15};
parameter YY15XX20={4'd15,4'd15,4'd15};
parameter YY15XX21={4'd15,4'd15,4'd15};
parameter YY15XX22={4'd15,4'd15,4'd15};
parameter YY15XX23={4'd15,4'd15,4'd15};
parameter YY15XX24={4'd15,4'd15,4'd14};
parameter YY15XX25={4'd10,4'd9,4'd9};
parameter YY15XX26={4'd15,4'd0,4'd0};
parameter YY15XX27={4'd15,4'd0,4'd0};
parameter YY15XX28={4'd15,4'd0,4'd0};
parameter YY16XX1={4'd15,4'd0,4'd0};
parameter YY16XX2={4'd5,4'd5,4'd4};
parameter YY16XX3={4'd9,4'd9,4'd8};
parameter YY16XX4={4'd13,4'd14,4'd13};
parameter YY16XX5={4'd14,4'd15,4'd15};
parameter YY16XX6={4'd15,4'd15,4'd15};
parameter YY16XX7={4'd15,4'd15,4'd15};
parameter YY16XX8={4'd15,4'd15,4'd15};
parameter YY16XX9={4'd15,4'd15,4'd15};
parameter YY16XX10={4'd15,4'd15,4'd15};
parameter YY16XX11={4'd15,4'd15,4'd15};
parameter YY16XX12={4'd15,4'd15,4'd15};
parameter YY16XX13={4'd15,4'd15,4'd15};
parameter YY16XX14={4'd15,4'd15,4'd15};
parameter YY16XX15={4'd15,4'd15,4'd15};
parameter YY16XX16={4'd15,4'd15,4'd15};
parameter YY16XX17={4'd15,4'd15,4'd15};
parameter YY16XX18={4'd15,4'd15,4'd15};
parameter YY16XX19={4'd15,4'd15,4'd15};
parameter YY16XX20={4'd15,4'd15,4'd15};
parameter YY16XX21={4'd15,4'd15,4'd15};
parameter YY16XX22={4'd15,4'd15,4'd15};
parameter YY16XX23={4'd15,4'd15,4'd15};
parameter YY16XX24={4'd14,4'd14,4'd14};
parameter YY16XX25={4'd9,4'd9,4'd8};
parameter YY16XX26={4'd15,4'd0,4'd0};
parameter YY16XX27={4'd15,4'd0,4'd0};
parameter YY16XX28={4'd15,4'd0,4'd0};
parameter YY17XX1={4'd15,4'd0,4'd0};
parameter YY17XX2={4'd4,4'd3,4'd3};
parameter YY17XX3={4'd8,4'd8,4'd7};
parameter YY17XX4={4'd13,4'd13,4'd13};
parameter YY17XX5={4'd14,4'd15,4'd15};
parameter YY17XX6={4'd15,4'd15,4'd15};
parameter YY17XX7={4'd15,4'd15,4'd15};
parameter YY17XX8={4'd15,4'd15,4'd15};
parameter YY17XX9={4'd15,4'd15,4'd15};
parameter YY17XX10={4'd15,4'd15,4'd15};
parameter YY17XX11={4'd15,4'd15,4'd15};
parameter YY17XX12={4'd15,4'd15,4'd15};
parameter YY17XX13={4'd15,4'd15,4'd15};
parameter YY17XX14={4'd15,4'd15,4'd15};
parameter YY17XX15={4'd15,4'd15,4'd15};
parameter YY17XX16={4'd15,4'd15,4'd15};
parameter YY17XX17={4'd15,4'd15,4'd15};
parameter YY17XX18={4'd15,4'd15,4'd15};
parameter YY17XX19={4'd15,4'd15,4'd15};
parameter YY17XX20={4'd15,4'd15,4'd15};
parameter YY17XX21={4'd15,4'd15,4'd15};
parameter YY17XX22={4'd15,4'd15,4'd15};
parameter YY17XX23={4'd15,4'd15,4'd15};
parameter YY17XX24={4'd14,4'd14,4'd14};
parameter YY17XX25={4'd8,4'd8,4'd8};
parameter YY17XX26={4'd15,4'd0,4'd0};
parameter YY17XX27={4'd15,4'd0,4'd0};
parameter YY17XX28={4'd15,4'd0,4'd0};
parameter YY18XX1={4'd15,4'd0,4'd0};
parameter YY18XX2={4'd5,4'd5,4'd4};
parameter YY18XX3={4'd9,4'd9,4'd8};
parameter YY18XX4={4'd13,4'd13,4'd13};
parameter YY18XX5={4'd14,4'd14,4'd14};
parameter YY18XX6={4'd15,4'd15,4'd15};
parameter YY18XX7={4'd15,4'd15,4'd15};
parameter YY18XX8={4'd15,4'd15,4'd15};
parameter YY18XX9={4'd15,4'd15,4'd15};
parameter YY18XX10={4'd15,4'd15,4'd15};
parameter YY18XX11={4'd15,4'd15,4'd15};
parameter YY18XX12={4'd15,4'd15,4'd15};
parameter YY18XX13={4'd15,4'd15,4'd15};
parameter YY18XX14={4'd15,4'd15,4'd15};
parameter YY18XX15={4'd15,4'd15,4'd15};
parameter YY18XX16={4'd15,4'd15,4'd15};
parameter YY18XX17={4'd15,4'd15,4'd15};
parameter YY18XX18={4'd15,4'd15,4'd15};
parameter YY18XX19={4'd15,4'd15,4'd15};
parameter YY18XX20={4'd15,4'd15,4'd15};
parameter YY18XX21={4'd15,4'd15,4'd15};
parameter YY18XX22={4'd15,4'd15,4'd15};
parameter YY18XX23={4'd15,4'd15,4'd15};
parameter YY18XX24={4'd14,4'd14,4'd14};
parameter YY18XX25={4'd8,4'd8,4'd8};
parameter YY18XX26={4'd15,4'd0,4'd0};
parameter YY18XX27={4'd15,4'd0,4'd0};
parameter YY18XX28={4'd15,4'd0,4'd0};
parameter YY19XX1={4'd6,4'd5,4'd3};
parameter YY19XX2={4'd9,4'd8,4'd7};
parameter YY19XX3={4'd11,4'd11,4'd11};
parameter YY19XX4={4'd14,4'd13,4'd13};
parameter YY19XX5={4'd14,4'd14,4'd14};
parameter YY19XX6={4'd15,4'd15,4'd15};
parameter YY19XX7={4'd15,4'd15,4'd15};
parameter YY19XX8={4'd15,4'd15,4'd15};
parameter YY19XX9={4'd15,4'd15,4'd15};
parameter YY19XX10={4'd15,4'd15,4'd15};
parameter YY19XX11={4'd15,4'd15,4'd15};
parameter YY19XX12={4'd15,4'd15,4'd15};
parameter YY19XX13={4'd15,4'd15,4'd15};
parameter YY19XX14={4'd15,4'd15,4'd15};
parameter YY19XX15={4'd15,4'd15,4'd15};
parameter YY19XX16={4'd15,4'd15,4'd15};
parameter YY19XX17={4'd15,4'd15,4'd15};
parameter YY19XX18={4'd15,4'd15,4'd15};
parameter YY19XX19={4'd15,4'd15,4'd15};
parameter YY19XX20={4'd15,4'd15,4'd15};
parameter YY19XX21={4'd15,4'd15,4'd15};
parameter YY19XX22={4'd15,4'd15,4'd15};
parameter YY19XX23={4'd15,4'd15,4'd15};
parameter YY19XX24={4'd13,4'd14,4'd13};
parameter YY19XX25={4'd8,4'd8,4'd7};
parameter YY19XX26={4'd15,4'd0,4'd0};
parameter YY19XX27={4'd15,4'd0,4'd0};
parameter YY19XX28={4'd15,4'd0,4'd0};
parameter YY20XX1={4'd7,4'd6,4'd4};
parameter YY20XX2={4'd11,4'd10,4'd9};
parameter YY20XX3={4'd14,4'd13,4'd13};
parameter YY20XX4={4'd15,4'd14,4'd14};
parameter YY20XX5={4'd14,4'd14,4'd14};
parameter YY20XX6={4'd15,4'd15,4'd15};
parameter YY20XX7={4'd15,4'd15,4'd15};
parameter YY20XX8={4'd15,4'd15,4'd15};
parameter YY20XX9={4'd15,4'd15,4'd15};
parameter YY20XX10={4'd15,4'd15,4'd15};
parameter YY20XX11={4'd15,4'd15,4'd15};
parameter YY20XX12={4'd15,4'd15,4'd15};
parameter YY20XX13={4'd15,4'd15,4'd15};
parameter YY20XX14={4'd15,4'd15,4'd15};
parameter YY20XX15={4'd15,4'd15,4'd15};
parameter YY20XX16={4'd15,4'd15,4'd15};
parameter YY20XX17={4'd15,4'd15,4'd15};
parameter YY20XX18={4'd15,4'd15,4'd15};
parameter YY20XX19={4'd15,4'd15,4'd15};
parameter YY20XX20={4'd15,4'd15,4'd15};
parameter YY20XX21={4'd15,4'd15,4'd15};
parameter YY20XX22={4'd15,4'd15,4'd15};
parameter YY20XX23={4'd15,4'd15,4'd15};
parameter YY20XX24={4'd13,4'd14,4'd13};
parameter YY20XX25={4'd7,4'd8,4'd7};
parameter YY20XX26={4'd15,4'd0,4'd0};
parameter YY20XX27={4'd15,4'd0,4'd0};
parameter YY20XX28={4'd15,4'd0,4'd0};
parameter YY21XX1={4'd9,4'd8,4'd6};
parameter YY21XX2={4'd12,4'd11,4'd10};
parameter YY21XX3={4'd15,4'd14,4'd14};
parameter YY21XX4={4'd15,4'd15,4'd15};
parameter YY21XX5={4'd15,4'd15,4'd15};
parameter YY21XX6={4'd15,4'd15,4'd15};
parameter YY21XX7={4'd15,4'd15,4'd15};
parameter YY21XX8={4'd15,4'd15,4'd15};
parameter YY21XX9={4'd15,4'd15,4'd15};
parameter YY21XX10={4'd15,4'd15,4'd15};
parameter YY21XX11={4'd15,4'd15,4'd15};
parameter YY21XX12={4'd15,4'd15,4'd15};
parameter YY21XX13={4'd15,4'd15,4'd15};
parameter YY21XX14={4'd15,4'd15,4'd15};
parameter YY21XX15={4'd15,4'd15,4'd15};
parameter YY21XX16={4'd15,4'd15,4'd15};
parameter YY21XX17={4'd15,4'd15,4'd15};
parameter YY21XX18={4'd15,4'd15,4'd15};
parameter YY21XX19={4'd15,4'd15,4'd15};
parameter YY21XX20={4'd15,4'd15,4'd15};
parameter YY21XX21={4'd15,4'd15,4'd15};
parameter YY21XX22={4'd15,4'd15,4'd15};
parameter YY21XX23={4'd15,4'd15,4'd15};
parameter YY21XX24={4'd12,4'd12,4'd12};
parameter YY21XX25={4'd7,4'd8,4'd7};
parameter YY21XX26={4'd15,4'd0,4'd0};
parameter YY21XX27={4'd15,4'd0,4'd0};
parameter YY21XX28={4'd15,4'd0,4'd0};
parameter YY22XX1={4'd10,4'd9,4'd8};
parameter YY22XX2={4'd13,4'd12,4'd11};
parameter YY22XX3={4'd15,4'd15,4'd14};
parameter YY22XX4={4'd15,4'd15,4'd15};
parameter YY22XX5={4'd15,4'd15,4'd15};
parameter YY22XX6={4'd15,4'd15,4'd15};
parameter YY22XX7={4'd15,4'd15,4'd15};
parameter YY22XX8={4'd15,4'd15,4'd15};
parameter YY22XX9={4'd15,4'd15,4'd15};
parameter YY22XX10={4'd15,4'd15,4'd15};
parameter YY22XX11={4'd15,4'd15,4'd15};
parameter YY22XX12={4'd15,4'd15,4'd15};
parameter YY22XX13={4'd15,4'd15,4'd15};
parameter YY22XX14={4'd15,4'd15,4'd15};
parameter YY22XX15={4'd15,4'd15,4'd15};
parameter YY22XX16={4'd15,4'd15,4'd15};
parameter YY22XX17={4'd15,4'd15,4'd15};
parameter YY22XX18={4'd15,4'd15,4'd15};
parameter YY22XX19={4'd15,4'd15,4'd15};
parameter YY22XX20={4'd15,4'd15,4'd15};
parameter YY22XX21={4'd15,4'd15,4'd15};
parameter YY22XX22={4'd15,4'd15,4'd15};
parameter YY22XX23={4'd14,4'd14,4'd14};
parameter YY22XX24={4'd12,4'd12,4'd12};
parameter YY22XX25={4'd9,4'd9,4'd9};
parameter YY22XX26={4'd7,4'd7,4'd7};
parameter YY22XX27={4'd5,4'd5,4'd5};
parameter YY22XX28={4'd15,4'd0,4'd0};
parameter YY23XX1={4'd11,4'd10,4'd9};
parameter YY23XX2={4'd13,4'd13,4'd12};
parameter YY23XX3={4'd15,4'd15,4'd15};
parameter YY23XX4={4'd15,4'd15,4'd15};
parameter YY23XX5={4'd15,4'd15,4'd15};
parameter YY23XX6={4'd15,4'd15,4'd15};
parameter YY23XX7={4'd15,4'd15,4'd15};
parameter YY23XX8={4'd15,4'd15,4'd15};
parameter YY23XX9={4'd15,4'd15,4'd15};
parameter YY23XX10={4'd15,4'd15,4'd15};
parameter YY23XX11={4'd15,4'd15,4'd15};
parameter YY23XX12={4'd15,4'd15,4'd15};
parameter YY23XX13={4'd15,4'd15,4'd15};
parameter YY23XX14={4'd15,4'd15,4'd15};
parameter YY23XX15={4'd15,4'd15,4'd15};
parameter YY23XX16={4'd15,4'd15,4'd15};
parameter YY23XX17={4'd15,4'd15,4'd15};
parameter YY23XX18={4'd15,4'd15,4'd15};
parameter YY23XX19={4'd15,4'd15,4'd15};
parameter YY23XX20={4'd15,4'd15,4'd15};
parameter YY23XX21={4'd15,4'd15,4'd15};
parameter YY23XX22={4'd14,4'd14,4'd14};
parameter YY23XX23={4'd11,4'd12,4'd11};
parameter YY23XX24={4'd11,4'd11,4'd11};
parameter YY23XX25={4'd11,4'd11,4'd11};
parameter YY23XX26={4'd12,4'd12,4'd12};
parameter YY23XX27={4'd11,4'd11,4'd11};
parameter YY23XX28={4'd8,4'd8,4'd7};
parameter YY24XX1={4'd9,4'd9,4'd8};
parameter YY24XX2={4'd11,4'd12,4'd11};
parameter YY24XX3={4'd14,4'd14,4'd14};
parameter YY24XX4={4'd15,4'd15,4'd15};
parameter YY24XX5={4'd15,4'd15,4'd15};
parameter YY24XX6={4'd15,4'd15,4'd15};
parameter YY24XX7={4'd15,4'd15,4'd15};
parameter YY24XX8={4'd15,4'd15,4'd15};
parameter YY24XX9={4'd15,4'd15,4'd15};
parameter YY24XX10={4'd15,4'd15,4'd15};
parameter YY24XX11={4'd15,4'd15,4'd15};
parameter YY24XX12={4'd15,4'd15,4'd15};
parameter YY24XX13={4'd15,4'd15,4'd15};
parameter YY24XX14={4'd15,4'd15,4'd15};
parameter YY24XX15={4'd15,4'd15,4'd15};
parameter YY24XX16={4'd15,4'd15,4'd15};
parameter YY24XX17={4'd15,4'd15,4'd15};
parameter YY24XX18={4'd15,4'd15,4'd15};
parameter YY24XX19={4'd15,4'd15,4'd15};
parameter YY24XX20={4'd15,4'd15,4'd15};
parameter YY24XX21={4'd15,4'd14,4'd15};
parameter YY24XX22={4'd14,4'd14,4'd14};
parameter YY24XX23={4'd14,4'd14,4'd14};
parameter YY24XX24={4'd13,4'd14,4'd14};
parameter YY24XX25={4'd14,4'd14,4'd14};
parameter YY24XX26={4'd15,4'd15,4'd15};
parameter YY24XX27={4'd14,4'd14,4'd14};
parameter YY24XX28={4'd10,4'd10,4'd9};
parameter YY25XX1={4'd6,4'd6,4'd6};
parameter YY25XX2={4'd8,4'd8,4'd8};
parameter YY25XX3={4'd11,4'd11,4'd11};
parameter YY25XX4={4'd13,4'd14,4'd14};
parameter YY25XX5={4'd14,4'd15,4'd15};
parameter YY25XX6={4'd15,4'd15,4'd15};
parameter YY25XX7={4'd15,4'd15,4'd15};
parameter YY25XX8={4'd15,4'd15,4'd15};
parameter YY25XX9={4'd15,4'd15,4'd15};
parameter YY25XX10={4'd15,4'd15,4'd15};
parameter YY25XX11={4'd15,4'd15,4'd15};
parameter YY25XX12={4'd15,4'd15,4'd15};
parameter YY25XX13={4'd15,4'd15,4'd15};
parameter YY25XX14={4'd15,4'd15,4'd15};
parameter YY25XX15={4'd15,4'd15,4'd15};
parameter YY25XX16={4'd15,4'd15,4'd15};
parameter YY25XX17={4'd15,4'd15,4'd15};
parameter YY25XX18={4'd15,4'd15,4'd15};
parameter YY25XX19={4'd15,4'd14,4'd15};
parameter YY25XX20={4'd15,4'd14,4'd14};
parameter YY25XX21={4'd15,4'd14,4'd15};
parameter YY25XX22={4'd14,4'd14,4'd14};
parameter YY25XX23={4'd15,4'd15,4'd15};
parameter YY25XX24={4'd15,4'd15,4'd15};
parameter YY25XX25={4'd15,4'd15,4'd15};
parameter YY25XX26={4'd15,4'd15,4'd15};
parameter YY25XX27={4'd12,4'd12,4'd11};
parameter YY25XX28={4'd7,4'd7,4'd6};
parameter YY26XX1={4'd3,4'd3,4'd3};
parameter YY26XX2={4'd5,4'd5,4'd5};
parameter YY26XX3={4'd7,4'd8,4'd8};
parameter YY26XX4={4'd11,4'd12,4'd12};
parameter YY26XX5={4'd12,4'd13,4'd14};
parameter YY26XX6={4'd14,4'd14,4'd15};
parameter YY26XX7={4'd14,4'd14,4'd15};
parameter YY26XX8={4'd15,4'd14,4'd15};
parameter YY26XX9={4'd15,4'd15,4'd15};
parameter YY26XX10={4'd15,4'd15,4'd15};
parameter YY26XX11={4'd15,4'd15,4'd15};
parameter YY26XX12={4'd15,4'd15,4'd15};
parameter YY26XX13={4'd15,4'd15,4'd15};
parameter YY26XX14={4'd15,4'd15,4'd15};
parameter YY26XX15={4'd15,4'd15,4'd15};
parameter YY26XX16={4'd15,4'd15,4'd15};
parameter YY26XX17={4'd15,4'd15,4'd15};
parameter YY26XX18={4'd14,4'd13,4'd14};
parameter YY26XX19={4'd13,4'd13,4'd13};
parameter YY26XX20={4'd14,4'd13,4'd14};
parameter YY26XX21={4'd15,4'd14,4'd15};
parameter YY26XX22={4'd15,4'd15,4'd15};
parameter YY26XX23={4'd15,4'd15,4'd15};
parameter YY26XX24={4'd15,4'd15,4'd15};
parameter YY26XX25={4'd15,4'd15,4'd15};
parameter YY26XX26={4'd11,4'd11,4'd11};
parameter YY26XX27={4'd7,4'd7,4'd6};
parameter YY26XX28={4'd3,4'd3,4'd3};
parameter YY27XX1={4'd15,4'd0,4'd0};
parameter YY27XX2={4'd2,4'd3,4'd3};
parameter YY27XX3={4'd4,4'd5,4'd5};
parameter YY27XX4={4'd7,4'd8,4'd8};
parameter YY27XX5={4'd9,4'd10,4'd10};
parameter YY27XX6={4'd12,4'd12,4'd13};
parameter YY27XX7={4'd13,4'd13,4'd13};
parameter YY27XX8={4'd13,4'd13,4'd14};
parameter YY27XX9={4'd14,4'd13,4'd14};
parameter YY27XX10={4'd14,4'd14,4'd14};
parameter YY27XX11={4'd14,4'd14,4'd15};
parameter YY27XX12={4'd15,4'd14,4'd15};
parameter YY27XX13={4'd15,4'd14,4'd15};
parameter YY27XX14={4'd15,4'd14,4'd15};
parameter YY27XX15={4'd15,4'd14,4'd15};
parameter YY27XX16={4'd14,4'd14,4'd14};
parameter YY27XX17={4'd13,4'd13,4'd13};
parameter YY27XX18={4'd12,4'd12,4'd12};
parameter YY27XX19={4'd12,4'd12,4'd12};
parameter YY27XX20={4'd14,4'd13,4'd14};
parameter YY27XX21={4'd15,4'd15,4'd15};
parameter YY27XX22={4'd15,4'd15,4'd15};
parameter YY27XX23={4'd15,4'd15,4'd15};
parameter YY27XX24={4'd15,4'd15,4'd15};
parameter YY27XX25={4'd11,4'd11,4'd11};
parameter YY27XX26={4'd7,4'd7,4'd7};
parameter YY27XX27={4'd3,4'd3,4'd3};
parameter YY27XX28={4'd15,4'd0,4'd0};
parameter YY28XX1={4'd15,4'd0,4'd0};
parameter YY28XX2={4'd15,4'd0,4'd0};
parameter YY28XX3={4'd2,4'd2,4'd2};
parameter YY28XX4={4'd4,4'd4,4'd5};
parameter YY28XX5={4'd6,4'd6,4'd7};
parameter YY28XX6={4'd9,4'd9,4'd10};
parameter YY28XX7={4'd11,4'd11,4'd12};
parameter YY28XX8={4'd12,4'd11,4'd12};
parameter YY28XX9={4'd12,4'd12,4'd12};
parameter YY28XX10={4'd12,4'd12,4'd12};
parameter YY28XX11={4'd13,4'd12,4'd13};
parameter YY28XX12={4'd13,4'd12,4'd13};
parameter YY28XX13={4'd13,4'd12,4'd13};
parameter YY28XX14={4'd13,4'd12,4'd13};
parameter YY28XX15={4'd13,4'd12,4'd13};
parameter YY28XX16={4'd12,4'd12,4'd12};
parameter YY28XX17={4'd11,4'd11,4'd11};
parameter YY28XX18={4'd11,4'd11,4'd11};
parameter YY28XX19={4'd12,4'd12,4'd12};
parameter YY28XX20={4'd15,4'd14,4'd15};
parameter YY28XX21={4'd15,4'd15,4'd15};
parameter YY28XX22={4'd15,4'd15,4'd15};
parameter YY28XX23={4'd14,4'd14,4'd14};
parameter YY28XX24={4'd11,4'd11,4'd11};
parameter YY28XX25={4'd6,4'd6,4'd6};
parameter YY28XX26={4'd2,4'd2,4'd2};
parameter YY28XX27={4'd15,4'd0,4'd0};
parameter YY28XX28={4'd15,4'd0,4'd0};
parameter YY29XX1={4'd15,4'd0,4'd0};
parameter YY29XX2={4'd15,4'd0,4'd0};
parameter YY29XX3={4'd15,4'd0,4'd0};
parameter YY29XX4={4'd15,4'd0,4'd0};
parameter YY29XX5={4'd4,4'd3,4'd3};
parameter YY29XX6={4'd5,4'd5,4'd5};
parameter YY29XX7={4'd8,4'd7,4'd8};
parameter YY29XX8={4'd9,4'd8,4'd8};
parameter YY29XX9={4'd9,4'd9,4'd9};
parameter YY29XX10={4'd9,4'd9,4'd9};
parameter YY29XX11={4'd9,4'd9,4'd9};
parameter YY29XX12={4'd9,4'd9,4'd10};
parameter YY29XX13={4'd10,4'd9,4'd10};
parameter YY29XX14={4'd9,4'd9,4'd9};
parameter YY29XX15={4'd8,4'd8,4'd8};
parameter YY29XX16={4'd9,4'd9,4'd9};
parameter YY29XX17={4'd10,4'd9,4'd10};
parameter YY29XX18={4'd11,4'd11,4'd11};
parameter YY29XX19={4'd13,4'd13,4'd14};
parameter YY29XX20={4'd15,4'd15,4'd15};
parameter YY29XX21={4'd15,4'd15,4'd15};
parameter YY29XX22={4'd13,4'd13,4'd13};
parameter YY29XX23={4'd8,4'd8,4'd8};
parameter YY29XX24={4'd5,4'd5,4'd4};
parameter YY29XX25={4'd1,4'd1,4'd1};
parameter YY29XX26={4'd15,4'd0,4'd0};
parameter YY29XX27={4'd15,4'd0,4'd0};
parameter YY29XX28={4'd15,4'd0,4'd0};
parameter YY30XX1={4'd15,4'd0,4'd0};
parameter YY30XX2={4'd15,4'd0,4'd0};
parameter YY30XX3={4'd15,4'd0,4'd0};
parameter YY30XX4={4'd15,4'd0,4'd0};
parameter YY30XX5={4'd15,4'd0,4'd0};
parameter YY30XX6={4'd3,4'd2,4'd2};
parameter YY30XX7={4'd4,4'd4,4'd4};
parameter YY30XX8={4'd5,4'd5,4'd5};
parameter YY30XX9={4'd6,4'd6,4'd6};
parameter YY30XX10={4'd7,4'd7,4'd7};
parameter YY30XX11={4'd7,4'd7,4'd7};
parameter YY30XX12={4'd6,4'd6,4'd6};
parameter YY30XX13={4'd6,4'd6,4'd6};
parameter YY30XX14={4'd7,4'd6,4'd7};
parameter YY30XX15={4'd7,4'd6,4'd7};
parameter YY30XX16={4'd7,4'd7,4'd7};
parameter YY30XX17={4'd9,4'd8,4'd9};
parameter YY30XX18={4'd11,4'd10,4'd11};
parameter YY30XX19={4'd13,4'd13,4'd13};
parameter YY30XX20={4'd14,4'd14,4'd14};
parameter YY30XX21={4'd11,4'd11,4'd11};
parameter YY30XX22={4'd7,4'd7,4'd7};
parameter YY30XX23={4'd5,4'd4,4'd4};
parameter YY30XX24={4'd3,4'd3,4'd2};
parameter YY30XX25={4'd15,4'd0,4'd0};
parameter YY30XX26={4'd15,4'd0,4'd0};
parameter YY30XX27={4'd15,4'd0,4'd0};
parameter YY30XX28={4'd15,4'd0,4'd0};
parameter YY31XX1={4'd15,4'd0,4'd0};
parameter YY31XX2={4'd15,4'd0,4'd0};
parameter YY31XX3={4'd15,4'd0,4'd0};
parameter YY31XX4={4'd15,4'd0,4'd0};
parameter YY31XX5={4'd15,4'd0,4'd0};
parameter YY31XX6={4'd15,4'd0,4'd0};
parameter YY31XX7={4'd15,4'd0,4'd0};
parameter YY31XX8={4'd3,4'd3,4'd3};
parameter YY31XX9={4'd5,4'd4,4'd4};
parameter YY31XX10={4'd6,4'd6,4'd6};
parameter YY31XX11={4'd5,4'd5,4'd5};
parameter YY31XX12={4'd5,4'd4,4'd4};
parameter YY31XX13={4'd5,4'd5,4'd5};
parameter YY31XX14={4'd6,4'd6,4'd6};
parameter YY31XX15={4'd7,4'd6,4'd7};
parameter YY31XX16={4'd8,4'd8,4'd8};
parameter YY31XX17={4'd9,4'd9,4'd9};
parameter YY31XX18={4'd11,4'd10,4'd11};
parameter YY31XX19={4'd12,4'd12,4'd12};
parameter YY31XX20={4'd11,4'd11,4'd11};
parameter YY31XX21={4'd7,4'd7,4'd7};
parameter YY31XX22={4'd3,4'd2,4'd3};
parameter YY31XX23={4'd2,4'd2,4'd2};
parameter YY31XX24={4'd15,4'd0,4'd0};
parameter YY31XX25={4'd15,4'd0,4'd0};
parameter YY31XX26={4'd15,4'd0,4'd0};
parameter YY31XX27={4'd15,4'd0,4'd0};
parameter YY31XX28={4'd15,4'd0,4'd0};
parameter YY32XX1={4'd15,4'd0,4'd0};
parameter YY32XX2={4'd15,4'd0,4'd0};
parameter YY32XX3={4'd15,4'd0,4'd0};
parameter YY32XX4={4'd15,4'd0,4'd0};
parameter YY32XX5={4'd15,4'd0,4'd0};
parameter YY32XX6={4'd15,4'd0,4'd0};
parameter YY32XX7={4'd15,4'd0,4'd0};
parameter YY32XX8={4'd15,4'd0,4'd0};
parameter YY32XX9={4'd15,4'd0,4'd0};
parameter YY32XX10={4'd15,4'd0,4'd0};
parameter YY32XX11={4'd15,4'd0,4'd0};
parameter YY32XX12={4'd15,4'd0,4'd0};
parameter YY32XX13={4'd15,4'd0,4'd0};
parameter YY32XX14={4'd5,4'd5,4'd5};
parameter YY32XX15={4'd8,4'd7,4'd7};
parameter YY32XX16={4'd10,4'd9,4'd9};
parameter YY32XX17={4'd11,4'd10,4'd10};
parameter YY32XX18={4'd10,4'd9,4'd10};
parameter YY32XX19={4'd8,4'd7,4'd8};
parameter YY32XX20={4'd6,4'd5,4'd6};
parameter YY32XX21={4'd4,4'd3,4'd4};
parameter YY32XX22={4'd2,4'd2,4'd2};
parameter YY32XX23={4'd15,4'd0,4'd0};
parameter YY32XX24={4'd15,4'd0,4'd0};
parameter YY32XX25={4'd15,4'd0,4'd0};
parameter YY32XX26={4'd15,4'd0,4'd0};
parameter YY32XX27={4'd15,4'd0,4'd0};
parameter YY32XX28={4'd15,4'd0,4'd0};
parameter YY33XX1={4'd15,4'd0,4'd0};
parameter YY33XX2={4'd15,4'd0,4'd0};
parameter YY33XX3={4'd15,4'd0,4'd0};
parameter YY33XX4={4'd15,4'd0,4'd0};
parameter YY33XX5={4'd15,4'd0,4'd0};
parameter YY33XX6={4'd15,4'd0,4'd0};
parameter YY33XX7={4'd15,4'd0,4'd0};
parameter YY33XX8={4'd15,4'd0,4'd0};
parameter YY33XX9={4'd15,4'd0,4'd0};
parameter YY33XX10={4'd15,4'd0,4'd0};
parameter YY33XX11={4'd15,4'd0,4'd0};
parameter YY33XX12={4'd15,4'd0,4'd0};
parameter YY33XX13={4'd15,4'd0,4'd0};
parameter YY33XX14={4'd4,4'd4,4'd3};
parameter YY33XX15={4'd7,4'd7,4'd6};
parameter YY33XX16={4'd8,4'd8,4'd8};
parameter YY33XX17={4'd8,4'd8,4'd8};
parameter YY33XX18={4'd6,4'd6,4'd6};
parameter YY33XX19={4'd3,4'd3,4'd3};
parameter YY33XX20={4'd2,4'd2,4'd2};
parameter YY33XX21={4'd2,4'd2,4'd2};
parameter YY33XX22={4'd15,4'd0,4'd0};
parameter YY33XX23={4'd15,4'd0,4'd0};
parameter YY33XX24={4'd15,4'd0,4'd0};
parameter YY33XX25={4'd15,4'd0,4'd0};
parameter YY33XX26={4'd15,4'd0,4'd0};
parameter YY33XX27={4'd15,4'd0,4'd0};
parameter YY33XX28={4'd15,4'd0,4'd0};
parameter YY34XX1={4'd15,4'd0,4'd0};
parameter YY34XX2={4'd15,4'd0,4'd0};
parameter YY34XX3={4'd15,4'd0,4'd0};
parameter YY34XX4={4'd15,4'd0,4'd0};
parameter YY34XX5={4'd15,4'd0,4'd0};
parameter YY34XX6={4'd15,4'd0,4'd0};
parameter YY34XX7={4'd15,4'd0,4'd0};
parameter YY34XX8={4'd15,4'd0,4'd0};
parameter YY34XX9={4'd15,4'd0,4'd0};
parameter YY34XX10={4'd15,4'd0,4'd0};
parameter YY34XX11={4'd15,4'd0,4'd0};
parameter YY34XX12={4'd15,4'd0,4'd0};
parameter YY34XX13={4'd15,4'd0,4'd0};
parameter YY34XX14={4'd3,4'd3,4'd2};
parameter YY34XX15={4'd5,4'd4,4'd4};
parameter YY34XX16={4'd5,4'd5,4'd4};
parameter YY34XX17={4'd4,4'd4,4'd4};
parameter YY34XX18={4'd3,4'd3,4'd3};
parameter YY34XX19={4'd2,4'd2,4'd2};
parameter YY34XX20={4'd15,4'd0,4'd0};
parameter YY34XX21={4'd15,4'd0,4'd0};
parameter YY34XX22={4'd15,4'd0,4'd0};
parameter YY34XX23={4'd15,4'd0,4'd0};
parameter YY34XX24={4'd15,4'd0,4'd0};
parameter YY34XX25={4'd15,4'd0,4'd0};
parameter YY34XX26={4'd15,4'd0,4'd0};
parameter YY34XX27={4'd15,4'd0,4'd0};
parameter YY34XX28={4'd15,4'd0,4'd0};
parameter YY35XX1={4'd15,4'd0,4'd0};
parameter YY35XX2={4'd15,4'd0,4'd0};
parameter YY35XX3={4'd15,4'd0,4'd0};
parameter YY35XX4={4'd15,4'd0,4'd0};
parameter YY35XX5={4'd15,4'd0,4'd0};
parameter YY35XX6={4'd15,4'd0,4'd0};
parameter YY35XX7={4'd15,4'd0,4'd0};
parameter YY35XX8={4'd15,4'd0,4'd0};
parameter YY35XX9={4'd15,4'd0,4'd0};
parameter YY35XX10={4'd15,4'd0,4'd0};
parameter YY35XX11={4'd15,4'd0,4'd0};
parameter YY35XX12={4'd15,4'd0,4'd0};
parameter YY35XX13={4'd15,4'd0,4'd0};
parameter YY35XX14={4'd15,4'd0,4'd0};
parameter YY35XX15={4'd3,4'd3,4'd2};
parameter YY35XX16={4'd3,4'd2,4'd2};
parameter YY35XX17={4'd2,4'd2,4'd2};
parameter YY35XX18={4'd2,4'd2,4'd1};
parameter YY35XX19={4'd15,4'd0,4'd0};
parameter YY35XX20={4'd15,4'd0,4'd0};
parameter YY35XX21={4'd15,4'd0,4'd0};
parameter YY35XX22={4'd15,4'd0,4'd0};
parameter YY35XX23={4'd15,4'd0,4'd0};
parameter YY35XX24={4'd15,4'd0,4'd0};
parameter YY35XX25={4'd15,4'd0,4'd0};
parameter YY35XX26={4'd15,4'd0,4'd0};
parameter YY35XX27={4'd15,4'd0,4'd0};
parameter YY35XX28={4'd15,4'd0,4'd0};

always@*
begin
case(YX)
Y0X0: RGB=YY0XX0;
Y0X1: RGB=YY0XX1;
Y0X2: RGB=YY0XX2;
Y0X3: RGB=YY0XX3;
Y0X4: RGB=YY0XX4;
Y0X5: RGB=YY0XX5;
Y0X6: RGB=YY0XX6;
Y0X7: RGB=YY0XX7;
Y0X8: RGB=YY0XX8;
Y0X9: RGB=YY0XX9;
Y0X10: RGB=YY0XX10;
Y0X11: RGB=YY0XX11;
Y0X12: RGB=YY0XX12;
Y0X13: RGB=YY0XX13;
Y0X14: RGB=YY0XX14;
Y0X15: RGB=YY0XX15;
Y0X16: RGB=YY0XX16;
Y0X17: RGB=YY0XX17;
Y0X18: RGB=YY0XX18;
Y0X19: RGB=YY0XX19;
Y0X20: RGB=YY0XX20;
Y0X21: RGB=YY0XX21;
Y0X22: RGB=YY0XX22;
Y0X23: RGB=YY0XX23;
Y0X24: RGB=YY0XX24;
Y0X25: RGB=YY0XX25;
Y0X26: RGB=YY0XX26;
Y0X27: RGB=YY0XX27;
Y0X28: RGB=YY0XX28;
Y1X1: RGB=YY1XX1;
Y1X2: RGB=YY1XX2;
Y1X3: RGB=YY1XX3;
Y1X4: RGB=YY1XX4;
Y1X5: RGB=YY1XX5;
Y1X6: RGB=YY1XX6;
Y1X7: RGB=YY1XX7;
Y1X8: RGB=YY1XX8;
Y1X9: RGB=YY1XX9;
Y1X10: RGB=YY1XX10;
Y1X11: RGB=YY1XX11;
Y1X12: RGB=YY1XX12;
Y1X13: RGB=YY1XX13;
Y1X14: RGB=YY1XX14;
Y1X15: RGB=YY1XX15;
Y1X16: RGB=YY1XX16;
Y1X17: RGB=YY1XX17;
Y1X18: RGB=YY1XX18;
Y1X19: RGB=YY1XX19;
Y1X20: RGB=YY1XX20;
Y1X21: RGB=YY1XX21;
Y1X22: RGB=YY1XX22;
Y1X23: RGB=YY1XX23;
Y1X24: RGB=YY1XX24;
Y1X25: RGB=YY1XX25;
Y1X26: RGB=YY1XX26;
Y1X27: RGB=YY1XX27;
Y1X28: RGB=YY1XX28;
Y2X1: RGB=YY2XX1;
Y2X2: RGB=YY2XX2;
Y2X3: RGB=YY2XX3;
Y2X4: RGB=YY2XX4;
Y2X5: RGB=YY2XX5;
Y2X6: RGB=YY2XX6;
Y2X7: RGB=YY2XX7;
Y2X8: RGB=YY2XX8;
Y2X9: RGB=YY2XX9;
Y2X10: RGB=YY2XX10;
Y2X11: RGB=YY2XX11;
Y2X12: RGB=YY2XX12;
Y2X13: RGB=YY2XX13;
Y2X14: RGB=YY2XX14;
Y2X15: RGB=YY2XX15;
Y2X16: RGB=YY2XX16;
Y2X17: RGB=YY2XX17;
Y2X18: RGB=YY2XX18;
Y2X19: RGB=YY2XX19;
Y2X20: RGB=YY2XX20;
Y2X21: RGB=YY2XX21;
Y2X22: RGB=YY2XX22;
Y2X23: RGB=YY2XX23;
Y2X24: RGB=YY2XX24;
Y2X25: RGB=YY2XX25;
Y2X26: RGB=YY2XX26;
Y2X27: RGB=YY2XX27;
Y2X28: RGB=YY2XX28;
Y3X1: RGB=YY3XX1;
Y3X2: RGB=YY3XX2;
Y3X3: RGB=YY3XX3;
Y3X4: RGB=YY3XX4;
Y3X5: RGB=YY3XX5;
Y3X6: RGB=YY3XX6;
Y3X7: RGB=YY3XX7;
Y3X8: RGB=YY3XX8;
Y3X9: RGB=YY3XX9;
Y3X10: RGB=YY3XX10;
Y3X11: RGB=YY3XX11;
Y3X12: RGB=YY3XX12;
Y3X13: RGB=YY3XX13;
Y3X14: RGB=YY3XX14;
Y3X15: RGB=YY3XX15;
Y3X16: RGB=YY3XX16;
Y3X17: RGB=YY3XX17;
Y3X18: RGB=YY3XX18;
Y3X19: RGB=YY3XX19;
Y3X20: RGB=YY3XX20;
Y3X21: RGB=YY3XX21;
Y3X22: RGB=YY3XX22;
Y3X23: RGB=YY3XX23;
Y3X24: RGB=YY3XX24;
Y3X25: RGB=YY3XX25;
Y3X26: RGB=YY3XX26;
Y3X27: RGB=YY3XX27;
Y3X28: RGB=YY3XX28;
Y4X1: RGB=YY4XX1;
Y4X2: RGB=YY4XX2;
Y4X3: RGB=YY4XX3;
Y4X4: RGB=YY4XX4;
Y4X5: RGB=YY4XX5;
Y4X6: RGB=YY4XX6;
Y4X7: RGB=YY4XX7;
Y4X8: RGB=YY4XX8;
Y4X9: RGB=YY4XX9;
Y4X10: RGB=YY4XX10;
Y4X11: RGB=YY4XX11;
Y4X12: RGB=YY4XX12;
Y4X13: RGB=YY4XX13;
Y4X14: RGB=YY4XX14;
Y4X15: RGB=YY4XX15;
Y4X16: RGB=YY4XX16;
Y4X17: RGB=YY4XX17;
Y4X18: RGB=YY4XX18;
Y4X19: RGB=YY4XX19;
Y4X20: RGB=YY4XX20;
Y4X21: RGB=YY4XX21;
Y4X22: RGB=YY4XX22;
Y4X23: RGB=YY4XX23;
Y4X24: RGB=YY4XX24;
Y4X25: RGB=YY4XX25;
Y4X26: RGB=YY4XX26;
Y4X27: RGB=YY4XX27;
Y4X28: RGB=YY4XX28;
Y5X1: RGB=YY5XX1;
Y5X2: RGB=YY5XX2;
Y5X3: RGB=YY5XX3;
Y5X4: RGB=YY5XX4;
Y5X5: RGB=YY5XX5;
Y5X6: RGB=YY5XX6;
Y5X7: RGB=YY5XX7;
Y5X8: RGB=YY5XX8;
Y5X9: RGB=YY5XX9;
Y5X10: RGB=YY5XX10;
Y5X11: RGB=YY5XX11;
Y5X12: RGB=YY5XX12;
Y5X13: RGB=YY5XX13;
Y5X14: RGB=YY5XX14;
Y5X15: RGB=YY5XX15;
Y5X16: RGB=YY5XX16;
Y5X17: RGB=YY5XX17;
Y5X18: RGB=YY5XX18;
Y5X19: RGB=YY5XX19;
Y5X20: RGB=YY5XX20;
Y5X21: RGB=YY5XX21;
Y5X22: RGB=YY5XX22;
Y5X23: RGB=YY5XX23;
Y5X24: RGB=YY5XX24;
Y5X25: RGB=YY5XX25;
Y5X26: RGB=YY5XX26;
Y5X27: RGB=YY5XX27;
Y5X28: RGB=YY5XX28;
Y6X1: RGB=YY6XX1;
Y6X2: RGB=YY6XX2;
Y6X3: RGB=YY6XX3;
Y6X4: RGB=YY6XX4;
Y6X5: RGB=YY6XX5;
Y6X6: RGB=YY6XX6;
Y6X7: RGB=YY6XX7;
Y6X8: RGB=YY6XX8;
Y6X9: RGB=YY6XX9;
Y6X10: RGB=YY6XX10;
Y6X11: RGB=YY6XX11;
Y6X12: RGB=YY6XX12;
Y6X13: RGB=YY6XX13;
Y6X14: RGB=YY6XX14;
Y6X15: RGB=YY6XX15;
Y6X16: RGB=YY6XX16;
Y6X17: RGB=YY6XX17;
Y6X18: RGB=YY6XX18;
Y6X19: RGB=YY6XX19;
Y6X20: RGB=YY6XX20;
Y6X21: RGB=YY6XX21;
Y6X22: RGB=YY6XX22;
Y6X23: RGB=YY6XX23;
Y6X24: RGB=YY6XX24;
Y6X25: RGB=YY6XX25;
Y6X26: RGB=YY6XX26;
Y6X27: RGB=YY6XX27;
Y6X28: RGB=YY6XX28;
Y7X1: RGB=YY7XX1;
Y7X2: RGB=YY7XX2;
Y7X3: RGB=YY7XX3;
Y7X4: RGB=YY7XX4;
Y7X5: RGB=YY7XX5;
Y7X6: RGB=YY7XX6;
Y7X7: RGB=YY7XX7;
Y7X8: RGB=YY7XX8;
Y7X9: RGB=YY7XX9;
Y7X10: RGB=YY7XX10;
Y7X11: RGB=YY7XX11;
Y7X12: RGB=YY7XX12;
Y7X13: RGB=YY7XX13;
Y7X14: RGB=YY7XX14;
Y7X15: RGB=YY7XX15;
Y7X16: RGB=YY7XX16;
Y7X17: RGB=YY7XX17;
Y7X18: RGB=YY7XX18;
Y7X19: RGB=YY7XX19;
Y7X20: RGB=YY7XX20;
Y7X21: RGB=YY7XX21;
Y7X22: RGB=YY7XX22;
Y7X23: RGB=YY7XX23;
Y7X24: RGB=YY7XX24;
Y7X25: RGB=YY7XX25;
Y7X26: RGB=YY7XX26;
Y7X27: RGB=YY7XX27;
Y7X28: RGB=YY7XX28;
Y8X1: RGB=YY8XX1;
Y8X2: RGB=YY8XX2;
Y8X3: RGB=YY8XX3;
Y8X4: RGB=YY8XX4;
Y8X5: RGB=YY8XX5;
Y8X6: RGB=YY8XX6;
Y8X7: RGB=YY8XX7;
Y8X8: RGB=YY8XX8;
Y8X9: RGB=YY8XX9;
Y8X10: RGB=YY8XX10;
Y8X11: RGB=YY8XX11;
Y8X12: RGB=YY8XX12;
Y8X13: RGB=YY8XX13;
Y8X14: RGB=YY8XX14;
Y8X15: RGB=YY8XX15;
Y8X16: RGB=YY8XX16;
Y8X17: RGB=YY8XX17;
Y8X18: RGB=YY8XX18;
Y8X19: RGB=YY8XX19;
Y8X20: RGB=YY8XX20;
Y8X21: RGB=YY8XX21;
Y8X22: RGB=YY8XX22;
Y8X23: RGB=YY8XX23;
Y8X24: RGB=YY8XX24;
Y8X25: RGB=YY8XX25;
Y8X26: RGB=YY8XX26;
Y8X27: RGB=YY8XX27;
Y8X28: RGB=YY8XX28;
Y9X1: RGB=YY9XX1;
Y9X2: RGB=YY9XX2;
Y9X3: RGB=YY9XX3;
Y9X4: RGB=YY9XX4;
Y9X5: RGB=YY9XX5;
Y9X6: RGB=YY9XX6;
Y9X7: RGB=YY9XX7;
Y9X8: RGB=YY9XX8;
Y9X9: RGB=YY9XX9;
Y9X10: RGB=YY9XX10;
Y9X11: RGB=YY9XX11;
Y9X12: RGB=YY9XX12;
Y9X13: RGB=YY9XX13;
Y9X14: RGB=YY9XX14;
Y9X15: RGB=YY9XX15;
Y9X16: RGB=YY9XX16;
Y9X17: RGB=YY9XX17;
Y9X18: RGB=YY9XX18;
Y9X19: RGB=YY9XX19;
Y9X20: RGB=YY9XX20;
Y9X21: RGB=YY9XX21;
Y9X22: RGB=YY9XX22;
Y9X23: RGB=YY9XX23;
Y9X24: RGB=YY9XX24;
Y9X25: RGB=YY9XX25;
Y9X26: RGB=YY9XX26;
Y9X27: RGB=YY9XX27;
Y9X28: RGB=YY9XX28;
Y10X1: RGB=YY10XX1;
Y10X2: RGB=YY10XX2;
Y10X3: RGB=YY10XX3;
Y10X4: RGB=YY10XX4;
Y10X5: RGB=YY10XX5;
Y10X6: RGB=YY10XX6;
Y10X7: RGB=YY10XX7;
Y10X8: RGB=YY10XX8;
Y10X9: RGB=YY10XX9;
Y10X10: RGB=YY10XX10;
Y10X11: RGB=YY10XX11;
Y10X12: RGB=YY10XX12;
Y10X13: RGB=YY10XX13;
Y10X14: RGB=YY10XX14;
Y10X15: RGB=YY10XX15;
Y10X16: RGB=YY10XX16;
Y10X17: RGB=YY10XX17;
Y10X18: RGB=YY10XX18;
Y10X19: RGB=YY10XX19;
Y10X20: RGB=YY10XX20;
Y10X21: RGB=YY10XX21;
Y10X22: RGB=YY10XX22;
Y10X23: RGB=YY10XX23;
Y10X24: RGB=YY10XX24;
Y10X25: RGB=YY10XX25;
Y10X26: RGB=YY10XX26;
Y10X27: RGB=YY10XX27;
Y10X28: RGB=YY10XX28;
Y11X1: RGB=YY11XX1;
Y11X2: RGB=YY11XX2;
Y11X3: RGB=YY11XX3;
Y11X4: RGB=YY11XX4;
Y11X5: RGB=YY11XX5;
Y11X6: RGB=YY11XX6;
Y11X7: RGB=YY11XX7;
Y11X8: RGB=YY11XX8;
Y11X9: RGB=YY11XX9;
Y11X10: RGB=YY11XX10;
Y11X11: RGB=YY11XX11;
Y11X12: RGB=YY11XX12;
Y11X13: RGB=YY11XX13;
Y11X14: RGB=YY11XX14;
Y11X15: RGB=YY11XX15;
Y11X16: RGB=YY11XX16;
Y11X17: RGB=YY11XX17;
Y11X18: RGB=YY11XX18;
Y11X19: RGB=YY11XX19;
Y11X20: RGB=YY11XX20;
Y11X21: RGB=YY11XX21;
Y11X22: RGB=YY11XX22;
Y11X23: RGB=YY11XX23;
Y11X24: RGB=YY11XX24;
Y11X25: RGB=YY11XX25;
Y11X26: RGB=YY11XX26;
Y11X27: RGB=YY11XX27;
Y11X28: RGB=YY11XX28;
Y12X1: RGB=YY12XX1;
Y12X2: RGB=YY12XX2;
Y12X3: RGB=YY12XX3;
Y12X4: RGB=YY12XX4;
Y12X5: RGB=YY12XX5;
Y12X6: RGB=YY12XX6;
Y12X7: RGB=YY12XX7;
Y12X8: RGB=YY12XX8;
Y12X9: RGB=YY12XX9;
Y12X10: RGB=YY12XX10;
Y12X11: RGB=YY12XX11;
Y12X12: RGB=YY12XX12;
Y12X13: RGB=YY12XX13;
Y12X14: RGB=YY12XX14;
Y12X15: RGB=YY12XX15;
Y12X16: RGB=YY12XX16;
Y12X17: RGB=YY12XX17;
Y12X18: RGB=YY12XX18;
Y12X19: RGB=YY12XX19;
Y12X20: RGB=YY12XX20;
Y12X21: RGB=YY12XX21;
Y12X22: RGB=YY12XX22;
Y12X23: RGB=YY12XX23;
Y12X24: RGB=YY12XX24;
Y12X25: RGB=YY12XX25;
Y12X26: RGB=YY12XX26;
Y12X27: RGB=YY12XX27;
Y12X28: RGB=YY12XX28;
Y13X1: RGB=YY13XX1;
Y13X2: RGB=YY13XX2;
Y13X3: RGB=YY13XX3;
Y13X4: RGB=YY13XX4;
Y13X5: RGB=YY13XX5;
Y13X6: RGB=YY13XX6;
Y13X7: RGB=YY13XX7;
Y13X8: RGB=YY13XX8;
Y13X9: RGB=YY13XX9;
Y13X10: RGB=YY13XX10;
Y13X11: RGB=YY13XX11;
Y13X12: RGB=YY13XX12;
Y13X13: RGB=YY13XX13;
Y13X14: RGB=YY13XX14;
Y13X15: RGB=YY13XX15;
Y13X16: RGB=YY13XX16;
Y13X17: RGB=YY13XX17;
Y13X18: RGB=YY13XX18;
Y13X19: RGB=YY13XX19;
Y13X20: RGB=YY13XX20;
Y13X21: RGB=YY13XX21;
Y13X22: RGB=YY13XX22;
Y13X23: RGB=YY13XX23;
Y13X24: RGB=YY13XX24;
Y13X25: RGB=YY13XX25;
Y13X26: RGB=YY13XX26;
Y13X27: RGB=YY13XX27;
Y13X28: RGB=YY13XX28;
Y14X1: RGB=YY14XX1;
Y14X2: RGB=YY14XX2;
Y14X3: RGB=YY14XX3;
Y14X4: RGB=YY14XX4;
Y14X5: RGB=YY14XX5;
Y14X6: RGB=YY14XX6;
Y14X7: RGB=YY14XX7;
Y14X8: RGB=YY14XX8;
Y14X9: RGB=YY14XX9;
Y14X10: RGB=YY14XX10;
Y14X11: RGB=YY14XX11;
Y14X12: RGB=YY14XX12;
Y14X13: RGB=YY14XX13;
Y14X14: RGB=YY14XX14;
Y14X15: RGB=YY14XX15;
Y14X16: RGB=YY14XX16;
Y14X17: RGB=YY14XX17;
Y14X18: RGB=YY14XX18;
Y14X19: RGB=YY14XX19;
Y14X20: RGB=YY14XX20;
Y14X21: RGB=YY14XX21;
Y14X22: RGB=YY14XX22;
Y14X23: RGB=YY14XX23;
Y14X24: RGB=YY14XX24;
Y14X25: RGB=YY14XX25;
Y14X26: RGB=YY14XX26;
Y14X27: RGB=YY14XX27;
Y14X28: RGB=YY14XX28;
Y15X1: RGB=YY15XX1;
Y15X2: RGB=YY15XX2;
Y15X3: RGB=YY15XX3;
Y15X4: RGB=YY15XX4;
Y15X5: RGB=YY15XX5;
Y15X6: RGB=YY15XX6;
Y15X7: RGB=YY15XX7;
Y15X8: RGB=YY15XX8;
Y15X9: RGB=YY15XX9;
Y15X10: RGB=YY15XX10;
Y15X11: RGB=YY15XX11;
Y15X12: RGB=YY15XX12;
Y15X13: RGB=YY15XX13;
Y15X14: RGB=YY15XX14;
Y15X15: RGB=YY15XX15;
Y15X16: RGB=YY15XX16;
Y15X17: RGB=YY15XX17;
Y15X18: RGB=YY15XX18;
Y15X19: RGB=YY15XX19;
Y15X20: RGB=YY15XX20;
Y15X21: RGB=YY15XX21;
Y15X22: RGB=YY15XX22;
Y15X23: RGB=YY15XX23;
Y15X24: RGB=YY15XX24;
Y15X25: RGB=YY15XX25;
Y15X26: RGB=YY15XX26;
Y15X27: RGB=YY15XX27;
Y15X28: RGB=YY15XX28;
Y16X1: RGB=YY16XX1;
Y16X2: RGB=YY16XX2;
Y16X3: RGB=YY16XX3;
Y16X4: RGB=YY16XX4;
Y16X5: RGB=YY16XX5;
Y16X6: RGB=YY16XX6;
Y16X7: RGB=YY16XX7;
Y16X8: RGB=YY16XX8;
Y16X9: RGB=YY16XX9;
Y16X10: RGB=YY16XX10;
Y16X11: RGB=YY16XX11;
Y16X12: RGB=YY16XX12;
Y16X13: RGB=YY16XX13;
Y16X14: RGB=YY16XX14;
Y16X15: RGB=YY16XX15;
Y16X16: RGB=YY16XX16;
Y16X17: RGB=YY16XX17;
Y16X18: RGB=YY16XX18;
Y16X19: RGB=YY16XX19;
Y16X20: RGB=YY16XX20;
Y16X21: RGB=YY16XX21;
Y16X22: RGB=YY16XX22;
Y16X23: RGB=YY16XX23;
Y16X24: RGB=YY16XX24;
Y16X25: RGB=YY16XX25;
Y16X26: RGB=YY16XX26;
Y16X27: RGB=YY16XX27;
Y16X28: RGB=YY16XX28;
Y17X1: RGB=YY17XX1;
Y17X2: RGB=YY17XX2;
Y17X3: RGB=YY17XX3;
Y17X4: RGB=YY17XX4;
Y17X5: RGB=YY17XX5;
Y17X6: RGB=YY17XX6;
Y17X7: RGB=YY17XX7;
Y17X8: RGB=YY17XX8;
Y17X9: RGB=YY17XX9;
Y17X10: RGB=YY17XX10;
Y17X11: RGB=YY17XX11;
Y17X12: RGB=YY17XX12;
Y17X13: RGB=YY17XX13;
Y17X14: RGB=YY17XX14;
Y17X15: RGB=YY17XX15;
Y17X16: RGB=YY17XX16;
Y17X17: RGB=YY17XX17;
Y17X18: RGB=YY17XX18;
Y17X19: RGB=YY17XX19;
Y17X20: RGB=YY17XX20;
Y17X21: RGB=YY17XX21;
Y17X22: RGB=YY17XX22;
Y17X23: RGB=YY17XX23;
Y17X24: RGB=YY17XX24;
Y17X25: RGB=YY17XX25;
Y17X26: RGB=YY17XX26;
Y17X27: RGB=YY17XX27;
Y17X28: RGB=YY17XX28;
Y18X1: RGB=YY18XX1;
Y18X2: RGB=YY18XX2;
Y18X3: RGB=YY18XX3;
Y18X4: RGB=YY18XX4;
Y18X5: RGB=YY18XX5;
Y18X6: RGB=YY18XX6;
Y18X7: RGB=YY18XX7;
Y18X8: RGB=YY18XX8;
Y18X9: RGB=YY18XX9;
Y18X10: RGB=YY18XX10;
Y18X11: RGB=YY18XX11;
Y18X12: RGB=YY18XX12;
Y18X13: RGB=YY18XX13;
Y18X14: RGB=YY18XX14;
Y18X15: RGB=YY18XX15;
Y18X16: RGB=YY18XX16;
Y18X17: RGB=YY18XX17;
Y18X18: RGB=YY18XX18;
Y18X19: RGB=YY18XX19;
Y18X20: RGB=YY18XX20;
Y18X21: RGB=YY18XX21;
Y18X22: RGB=YY18XX22;
Y18X23: RGB=YY18XX23;
Y18X24: RGB=YY18XX24;
Y18X25: RGB=YY18XX25;
Y18X26: RGB=YY18XX26;
Y18X27: RGB=YY18XX27;
Y18X28: RGB=YY18XX28;
Y19X1: RGB=YY19XX1;
Y19X2: RGB=YY19XX2;
Y19X3: RGB=YY19XX3;
Y19X4: RGB=YY19XX4;
Y19X5: RGB=YY19XX5;
Y19X6: RGB=YY19XX6;
Y19X7: RGB=YY19XX7;
Y19X8: RGB=YY19XX8;
Y19X9: RGB=YY19XX9;
Y19X10: RGB=YY19XX10;
Y19X11: RGB=YY19XX11;
Y19X12: RGB=YY19XX12;
Y19X13: RGB=YY19XX13;
Y19X14: RGB=YY19XX14;
Y19X15: RGB=YY19XX15;
Y19X16: RGB=YY19XX16;
Y19X17: RGB=YY19XX17;
Y19X18: RGB=YY19XX18;
Y19X19: RGB=YY19XX19;
Y19X20: RGB=YY19XX20;
Y19X21: RGB=YY19XX21;
Y19X22: RGB=YY19XX22;
Y19X23: RGB=YY19XX23;
Y19X24: RGB=YY19XX24;
Y19X25: RGB=YY19XX25;
Y19X26: RGB=YY19XX26;
Y19X27: RGB=YY19XX27;
Y19X28: RGB=YY19XX28;
Y20X1: RGB=YY20XX1;
Y20X2: RGB=YY20XX2;
Y20X3: RGB=YY20XX3;
Y20X4: RGB=YY20XX4;
Y20X5: RGB=YY20XX5;
Y20X6: RGB=YY20XX6;
Y20X7: RGB=YY20XX7;
Y20X8: RGB=YY20XX8;
Y20X9: RGB=YY20XX9;
Y20X10: RGB=YY20XX10;
Y20X11: RGB=YY20XX11;
Y20X12: RGB=YY20XX12;
Y20X13: RGB=YY20XX13;
Y20X14: RGB=YY20XX14;
Y20X15: RGB=YY20XX15;
Y20X16: RGB=YY20XX16;
Y20X17: RGB=YY20XX17;
Y20X18: RGB=YY20XX18;
Y20X19: RGB=YY20XX19;
Y20X20: RGB=YY20XX20;
Y20X21: RGB=YY20XX21;
Y20X22: RGB=YY20XX22;
Y20X23: RGB=YY20XX23;
Y20X24: RGB=YY20XX24;
Y20X25: RGB=YY20XX25;
Y20X26: RGB=YY20XX26;
Y20X27: RGB=YY20XX27;
Y20X28: RGB=YY20XX28;
Y21X1: RGB=YY21XX1;
Y21X2: RGB=YY21XX2;
Y21X3: RGB=YY21XX3;
Y21X4: RGB=YY21XX4;
Y21X5: RGB=YY21XX5;
Y21X6: RGB=YY21XX6;
Y21X7: RGB=YY21XX7;
Y21X8: RGB=YY21XX8;
Y21X9: RGB=YY21XX9;
Y21X10: RGB=YY21XX10;
Y21X11: RGB=YY21XX11;
Y21X12: RGB=YY21XX12;
Y21X13: RGB=YY21XX13;
Y21X14: RGB=YY21XX14;
Y21X15: RGB=YY21XX15;
Y21X16: RGB=YY21XX16;
Y21X17: RGB=YY21XX17;
Y21X18: RGB=YY21XX18;
Y21X19: RGB=YY21XX19;
Y21X20: RGB=YY21XX20;
Y21X21: RGB=YY21XX21;
Y21X22: RGB=YY21XX22;
Y21X23: RGB=YY21XX23;
Y21X24: RGB=YY21XX24;
Y21X25: RGB=YY21XX25;
Y21X26: RGB=YY21XX26;
Y21X27: RGB=YY21XX27;
Y21X28: RGB=YY21XX28;
Y22X1: RGB=YY22XX1;
Y22X2: RGB=YY22XX2;
Y22X3: RGB=YY22XX3;
Y22X4: RGB=YY22XX4;
Y22X5: RGB=YY22XX5;
Y22X6: RGB=YY22XX6;
Y22X7: RGB=YY22XX7;
Y22X8: RGB=YY22XX8;
Y22X9: RGB=YY22XX9;
Y22X10: RGB=YY22XX10;
Y22X11: RGB=YY22XX11;
Y22X12: RGB=YY22XX12;
Y22X13: RGB=YY22XX13;
Y22X14: RGB=YY22XX14;
Y22X15: RGB=YY22XX15;
Y22X16: RGB=YY22XX16;
Y22X17: RGB=YY22XX17;
Y22X18: RGB=YY22XX18;
Y22X19: RGB=YY22XX19;
Y22X20: RGB=YY22XX20;
Y22X21: RGB=YY22XX21;
Y22X22: RGB=YY22XX22;
Y22X23: RGB=YY22XX23;
Y22X24: RGB=YY22XX24;
Y22X25: RGB=YY22XX25;
Y22X26: RGB=YY22XX26;
Y22X27: RGB=YY22XX27;
Y22X28: RGB=YY22XX28;
Y23X1: RGB=YY23XX1;
Y23X2: RGB=YY23XX2;
Y23X3: RGB=YY23XX3;
Y23X4: RGB=YY23XX4;
Y23X5: RGB=YY23XX5;
Y23X6: RGB=YY23XX6;
Y23X7: RGB=YY23XX7;
Y23X8: RGB=YY23XX8;
Y23X9: RGB=YY23XX9;
Y23X10: RGB=YY23XX10;
Y23X11: RGB=YY23XX11;
Y23X12: RGB=YY23XX12;
Y23X13: RGB=YY23XX13;
Y23X14: RGB=YY23XX14;
Y23X15: RGB=YY23XX15;
Y23X16: RGB=YY23XX16;
Y23X17: RGB=YY23XX17;
Y23X18: RGB=YY23XX18;
Y23X19: RGB=YY23XX19;
Y23X20: RGB=YY23XX20;
Y23X21: RGB=YY23XX21;
Y23X22: RGB=YY23XX22;
Y23X23: RGB=YY23XX23;
Y23X24: RGB=YY23XX24;
Y23X25: RGB=YY23XX25;
Y23X26: RGB=YY23XX26;
Y23X27: RGB=YY23XX27;
Y23X28: RGB=YY23XX28;
Y24X1: RGB=YY24XX1;
Y24X2: RGB=YY24XX2;
Y24X3: RGB=YY24XX3;
Y24X4: RGB=YY24XX4;
Y24X5: RGB=YY24XX5;
Y24X6: RGB=YY24XX6;
Y24X7: RGB=YY24XX7;
Y24X8: RGB=YY24XX8;
Y24X9: RGB=YY24XX9;
Y24X10: RGB=YY24XX10;
Y24X11: RGB=YY24XX11;
Y24X12: RGB=YY24XX12;
Y24X13: RGB=YY24XX13;
Y24X14: RGB=YY24XX14;
Y24X15: RGB=YY24XX15;
Y24X16: RGB=YY24XX16;
Y24X17: RGB=YY24XX17;
Y24X18: RGB=YY24XX18;
Y24X19: RGB=YY24XX19;
Y24X20: RGB=YY24XX20;
Y24X21: RGB=YY24XX21;
Y24X22: RGB=YY24XX22;
Y24X23: RGB=YY24XX23;
Y24X24: RGB=YY24XX24;
Y24X25: RGB=YY24XX25;
Y24X26: RGB=YY24XX26;
Y24X27: RGB=YY24XX27;
Y24X28: RGB=YY24XX28;
Y25X1: RGB=YY25XX1;
Y25X2: RGB=YY25XX2;
Y25X3: RGB=YY25XX3;
Y25X4: RGB=YY25XX4;
Y25X5: RGB=YY25XX5;
Y25X6: RGB=YY25XX6;
Y25X7: RGB=YY25XX7;
Y25X8: RGB=YY25XX8;
Y25X9: RGB=YY25XX9;
Y25X10: RGB=YY25XX10;
Y25X11: RGB=YY25XX11;
Y25X12: RGB=YY25XX12;
Y25X13: RGB=YY25XX13;
Y25X14: RGB=YY25XX14;
Y25X15: RGB=YY25XX15;
Y25X16: RGB=YY25XX16;
Y25X17: RGB=YY25XX17;
Y25X18: RGB=YY25XX18;
Y25X19: RGB=YY25XX19;
Y25X20: RGB=YY25XX20;
Y25X21: RGB=YY25XX21;
Y25X22: RGB=YY25XX22;
Y25X23: RGB=YY25XX23;
Y25X24: RGB=YY25XX24;
Y25X25: RGB=YY25XX25;
Y25X26: RGB=YY25XX26;
Y25X27: RGB=YY25XX27;
Y25X28: RGB=YY25XX28;
Y26X1: RGB=YY26XX1;
Y26X2: RGB=YY26XX2;
Y26X3: RGB=YY26XX3;
Y26X4: RGB=YY26XX4;
Y26X5: RGB=YY26XX5;
Y26X6: RGB=YY26XX6;
Y26X7: RGB=YY26XX7;
Y26X8: RGB=YY26XX8;
Y26X9: RGB=YY26XX9;
Y26X10: RGB=YY26XX10;
Y26X11: RGB=YY26XX11;
Y26X12: RGB=YY26XX12;
Y26X13: RGB=YY26XX13;
Y26X14: RGB=YY26XX14;
Y26X15: RGB=YY26XX15;
Y26X16: RGB=YY26XX16;
Y26X17: RGB=YY26XX17;
Y26X18: RGB=YY26XX18;
Y26X19: RGB=YY26XX19;
Y26X20: RGB=YY26XX20;
Y26X21: RGB=YY26XX21;
Y26X22: RGB=YY26XX22;
Y26X23: RGB=YY26XX23;
Y26X24: RGB=YY26XX24;
Y26X25: RGB=YY26XX25;
Y26X26: RGB=YY26XX26;
Y26X27: RGB=YY26XX27;
Y26X28: RGB=YY26XX28;
Y27X1: RGB=YY27XX1;
Y27X2: RGB=YY27XX2;
Y27X3: RGB=YY27XX3;
Y27X4: RGB=YY27XX4;
Y27X5: RGB=YY27XX5;
Y27X6: RGB=YY27XX6;
Y27X7: RGB=YY27XX7;
Y27X8: RGB=YY27XX8;
Y27X9: RGB=YY27XX9;
Y27X10: RGB=YY27XX10;
Y27X11: RGB=YY27XX11;
Y27X12: RGB=YY27XX12;
Y27X13: RGB=YY27XX13;
Y27X14: RGB=YY27XX14;
Y27X15: RGB=YY27XX15;
Y27X16: RGB=YY27XX16;
Y27X17: RGB=YY27XX17;
Y27X18: RGB=YY27XX18;
Y27X19: RGB=YY27XX19;
Y27X20: RGB=YY27XX20;
Y27X21: RGB=YY27XX21;
Y27X22: RGB=YY27XX22;
Y27X23: RGB=YY27XX23;
Y27X24: RGB=YY27XX24;
Y27X25: RGB=YY27XX25;
Y27X26: RGB=YY27XX26;
Y27X27: RGB=YY27XX27;
Y27X28: RGB=YY27XX28;
Y28X1: RGB=YY28XX1;
Y28X2: RGB=YY28XX2;
Y28X3: RGB=YY28XX3;
Y28X4: RGB=YY28XX4;
Y28X5: RGB=YY28XX5;
Y28X6: RGB=YY28XX6;
Y28X7: RGB=YY28XX7;
Y28X8: RGB=YY28XX8;
Y28X9: RGB=YY28XX9;
Y28X10: RGB=YY28XX10;
Y28X11: RGB=YY28XX11;
Y28X12: RGB=YY28XX12;
Y28X13: RGB=YY28XX13;
Y28X14: RGB=YY28XX14;
Y28X15: RGB=YY28XX15;
Y28X16: RGB=YY28XX16;
Y28X17: RGB=YY28XX17;
Y28X18: RGB=YY28XX18;
Y28X19: RGB=YY28XX19;
Y28X20: RGB=YY28XX20;
Y28X21: RGB=YY28XX21;
Y28X22: RGB=YY28XX22;
Y28X23: RGB=YY28XX23;
Y28X24: RGB=YY28XX24;
Y28X25: RGB=YY28XX25;
Y28X26: RGB=YY28XX26;
Y28X27: RGB=YY28XX27;
Y28X28: RGB=YY28XX28;
Y29X1: RGB=YY29XX1;
Y29X2: RGB=YY29XX2;
Y29X3: RGB=YY29XX3;
Y29X4: RGB=YY29XX4;
Y29X5: RGB=YY29XX5;
Y29X6: RGB=YY29XX6;
Y29X7: RGB=YY29XX7;
Y29X8: RGB=YY29XX8;
Y29X9: RGB=YY29XX9;
Y29X10: RGB=YY29XX10;
Y29X11: RGB=YY29XX11;
Y29X12: RGB=YY29XX12;
Y29X13: RGB=YY29XX13;
Y29X14: RGB=YY29XX14;
Y29X15: RGB=YY29XX15;
Y29X16: RGB=YY29XX16;
Y29X17: RGB=YY29XX17;
Y29X18: RGB=YY29XX18;
Y29X19: RGB=YY29XX19;
Y29X20: RGB=YY29XX20;
Y29X21: RGB=YY29XX21;
Y29X22: RGB=YY29XX22;
Y29X23: RGB=YY29XX23;
Y29X24: RGB=YY29XX24;
Y29X25: RGB=YY29XX25;
Y29X26: RGB=YY29XX26;
Y29X27: RGB=YY29XX27;
Y29X28: RGB=YY29XX28;
Y30X1: RGB=YY30XX1;
Y30X2: RGB=YY30XX2;
Y30X3: RGB=YY30XX3;
Y30X4: RGB=YY30XX4;
Y30X5: RGB=YY30XX5;
Y30X6: RGB=YY30XX6;
Y30X7: RGB=YY30XX7;
Y30X8: RGB=YY30XX8;
Y30X9: RGB=YY30XX9;
Y30X10: RGB=YY30XX10;
Y30X11: RGB=YY30XX11;
Y30X12: RGB=YY30XX12;
Y30X13: RGB=YY30XX13;
Y30X14: RGB=YY30XX14;
Y30X15: RGB=YY30XX15;
Y30X16: RGB=YY30XX16;
Y30X17: RGB=YY30XX17;
Y30X18: RGB=YY30XX18;
Y30X19: RGB=YY30XX19;
Y30X20: RGB=YY30XX20;
Y30X21: RGB=YY30XX21;
Y30X22: RGB=YY30XX22;
Y30X23: RGB=YY30XX23;
Y30X24: RGB=YY30XX24;
Y30X25: RGB=YY30XX25;
Y30X26: RGB=YY30XX26;
Y30X27: RGB=YY30XX27;
Y30X28: RGB=YY30XX28;
Y31X1: RGB=YY31XX1;
Y31X2: RGB=YY31XX2;
Y31X3: RGB=YY31XX3;
Y31X4: RGB=YY31XX4;
Y31X5: RGB=YY31XX5;
Y31X6: RGB=YY31XX6;
Y31X7: RGB=YY31XX7;
Y31X8: RGB=YY31XX8;
Y31X9: RGB=YY31XX9;
Y31X10: RGB=YY31XX10;
Y31X11: RGB=YY31XX11;
Y31X12: RGB=YY31XX12;
Y31X13: RGB=YY31XX13;
Y31X14: RGB=YY31XX14;
Y31X15: RGB=YY31XX15;
Y31X16: RGB=YY31XX16;
Y31X17: RGB=YY31XX17;
Y31X18: RGB=YY31XX18;
Y31X19: RGB=YY31XX19;
Y31X20: RGB=YY31XX20;
Y31X21: RGB=YY31XX21;
Y31X22: RGB=YY31XX22;
Y31X23: RGB=YY31XX23;
Y31X24: RGB=YY31XX24;
Y31X25: RGB=YY31XX25;
Y31X26: RGB=YY31XX26;
Y31X27: RGB=YY31XX27;
Y31X28: RGB=YY31XX28;
Y32X1: RGB=YY32XX1;
Y32X2: RGB=YY32XX2;
Y32X3: RGB=YY32XX3;
Y32X4: RGB=YY32XX4;
Y32X5: RGB=YY32XX5;
Y32X6: RGB=YY32XX6;
Y32X7: RGB=YY32XX7;
Y32X8: RGB=YY32XX8;
Y32X9: RGB=YY32XX9;
Y32X10: RGB=YY32XX10;
Y32X11: RGB=YY32XX11;
Y32X12: RGB=YY32XX12;
Y32X13: RGB=YY32XX13;
Y32X14: RGB=YY32XX14;
Y32X15: RGB=YY32XX15;
Y32X16: RGB=YY32XX16;
Y32X17: RGB=YY32XX17;
Y32X18: RGB=YY32XX18;
Y32X19: RGB=YY32XX19;
Y32X20: RGB=YY32XX20;
Y32X21: RGB=YY32XX21;
Y32X22: RGB=YY32XX22;
Y32X23: RGB=YY32XX23;
Y32X24: RGB=YY32XX24;
Y32X25: RGB=YY32XX25;
Y32X26: RGB=YY32XX26;
Y32X27: RGB=YY32XX27;
Y32X28: RGB=YY32XX28;
Y33X1: RGB=YY33XX1;
Y33X2: RGB=YY33XX2;
Y33X3: RGB=YY33XX3;
Y33X4: RGB=YY33XX4;
Y33X5: RGB=YY33XX5;
Y33X6: RGB=YY33XX6;
Y33X7: RGB=YY33XX7;
Y33X8: RGB=YY33XX8;
Y33X9: RGB=YY33XX9;
Y33X10: RGB=YY33XX10;
Y33X11: RGB=YY33XX11;
Y33X12: RGB=YY33XX12;
Y33X13: RGB=YY33XX13;
Y33X14: RGB=YY33XX14;
Y33X15: RGB=YY33XX15;
Y33X16: RGB=YY33XX16;
Y33X17: RGB=YY33XX17;
Y33X18: RGB=YY33XX18;
Y33X19: RGB=YY33XX19;
Y33X20: RGB=YY33XX20;
Y33X21: RGB=YY33XX21;
Y33X22: RGB=YY33XX22;
Y33X23: RGB=YY33XX23;
Y33X24: RGB=YY33XX24;
Y33X25: RGB=YY33XX25;
Y33X26: RGB=YY33XX26;
Y33X27: RGB=YY33XX27;
Y33X28: RGB=YY33XX28;
Y34X1: RGB=YY34XX1;
Y34X2: RGB=YY34XX2;
Y34X3: RGB=YY34XX3;
Y34X4: RGB=YY34XX4;
Y34X5: RGB=YY34XX5;
Y34X6: RGB=YY34XX6;
Y34X7: RGB=YY34XX7;
Y34X8: RGB=YY34XX8;
Y34X9: RGB=YY34XX9;
Y34X10: RGB=YY34XX10;
Y34X11: RGB=YY34XX11;
Y34X12: RGB=YY34XX12;
Y34X13: RGB=YY34XX13;
Y34X14: RGB=YY34XX14;
Y34X15: RGB=YY34XX15;
Y34X16: RGB=YY34XX16;
Y34X17: RGB=YY34XX17;
Y34X18: RGB=YY34XX18;
Y34X19: RGB=YY34XX19;
Y34X20: RGB=YY34XX20;
Y34X21: RGB=YY34XX21;
Y34X22: RGB=YY34XX22;
Y34X23: RGB=YY34XX23;
Y34X24: RGB=YY34XX24;
Y34X25: RGB=YY34XX25;
Y34X26: RGB=YY34XX26;
Y34X27: RGB=YY34XX27;
Y34X28: RGB=YY34XX28;
Y35X1: RGB=YY35XX1;
Y35X2: RGB=YY35XX2;
Y35X3: RGB=YY35XX3;
Y35X4: RGB=YY35XX4;
Y35X5: RGB=YY35XX5;
Y35X6: RGB=YY35XX6;
Y35X7: RGB=YY35XX7;
Y35X8: RGB=YY35XX8;
Y35X9: RGB=YY35XX9;
Y35X10: RGB=YY35XX10;
Y35X11: RGB=YY35XX11;
Y35X12: RGB=YY35XX12;
Y35X13: RGB=YY35XX13;
Y35X14: RGB=YY35XX14;
Y35X15: RGB=YY35XX15;
Y35X16: RGB=YY35XX16;
Y35X17: RGB=YY35XX17;
Y35X18: RGB=YY35XX18;
Y35X19: RGB=YY35XX19;
Y35X20: RGB=YY35XX20;
Y35X21: RGB=YY35XX21;
Y35X22: RGB=YY35XX22;
Y35X23: RGB=YY35XX23;
Y35X24: RGB=YY35XX24;
Y35X25: RGB=YY35XX25;
Y35X26: RGB=YY35XX26;
Y35X27: RGB=YY35XX27;
Y35X28: RGB=YY35XX28;

default: RGB=12'd0;
endcase
end
endmodule